library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom1 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"d4efc287",
    12 => x"86c0c64e",
    13 => x"49d4efc2",
    14 => x"48e0dcc2",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087d6db",
    19 => x"1e87fc98",
    20 => x"1e731e72",
    21 => x"02114812",
    22 => x"c34b87ca",
    23 => x"739b98df",
    24 => x"87f00288",
    25 => x"4a264b26",
    26 => x"731e4f26",
    27 => x"c11e721e",
    28 => x"87ca048b",
    29 => x"02114812",
    30 => x"028887c4",
    31 => x"4a2687f1",
    32 => x"4f264b26",
    33 => x"731e741e",
    34 => x"c11e721e",
    35 => x"87d0048b",
    36 => x"02114812",
    37 => x"c34c87ca",
    38 => x"749c98df",
    39 => x"87eb0288",
    40 => x"4b264a26",
    41 => x"4f264c26",
    42 => x"8148731e",
    43 => x"c502a973",
    44 => x"05531287",
    45 => x"4f2687f6",
    46 => x"4a66c41e",
    47 => x"51124871",
    48 => x"2687fb05",
    49 => x"48111e4f",
    50 => x"7808d4ff",
    51 => x"c14866c4",
    52 => x"58a6c888",
    53 => x"ed059870",
    54 => x"1e4f2687",
    55 => x"c348d4ff",
    56 => x"516878ff",
    57 => x"c14866c4",
    58 => x"58a6c888",
    59 => x"eb059870",
    60 => x"1e4f2687",
    61 => x"d4ff1e73",
    62 => x"7bffc34b",
    63 => x"ffc34a6b",
    64 => x"c8496b7b",
    65 => x"c3b17232",
    66 => x"4a6b7bff",
    67 => x"b27131c8",
    68 => x"6b7bffc3",
    69 => x"7232c849",
    70 => x"c44871b1",
    71 => x"264d2687",
    72 => x"264b264c",
    73 => x"5b5e0e4f",
    74 => x"710e5d5c",
    75 => x"4cd4ff4a",
    76 => x"ffc34972",
    77 => x"c27c7199",
    78 => x"05bfe0dc",
    79 => x"66d087c8",
    80 => x"d430c948",
    81 => x"66d058a6",
    82 => x"c329d849",
    83 => x"7c7199ff",
    84 => x"d04966d0",
    85 => x"99ffc329",
    86 => x"66d07c71",
    87 => x"c329c849",
    88 => x"7c7199ff",
    89 => x"c34966d0",
    90 => x"7c7199ff",
    91 => x"29d04972",
    92 => x"7199ffc3",
    93 => x"c94b6c7c",
    94 => x"c34dfff0",
    95 => x"d005abff",
    96 => x"7cffc387",
    97 => x"8dc14b6c",
    98 => x"c387c602",
    99 => x"f002abff",
   100 => x"fe487387",
   101 => x"c01e87c7",
   102 => x"48d4ff49",
   103 => x"c178ffc3",
   104 => x"b7c8c381",
   105 => x"87f104a9",
   106 => x"731e4f26",
   107 => x"c487e71e",
   108 => x"c04bdff8",
   109 => x"f0ffc01e",
   110 => x"fd49f7c1",
   111 => x"86c487e7",
   112 => x"c005a8c1",
   113 => x"d4ff87ea",
   114 => x"78ffc348",
   115 => x"c0c0c0c1",
   116 => x"c01ec0c0",
   117 => x"e9c1f0e1",
   118 => x"87c9fd49",
   119 => x"987086c4",
   120 => x"ff87ca05",
   121 => x"ffc348d4",
   122 => x"cb48c178",
   123 => x"87e6fe87",
   124 => x"fe058bc1",
   125 => x"48c087fd",
   126 => x"1e87e6fc",
   127 => x"d4ff1e73",
   128 => x"78ffc348",
   129 => x"1ec04bd3",
   130 => x"c1f0ffc0",
   131 => x"d4fc49c1",
   132 => x"7086c487",
   133 => x"87ca0598",
   134 => x"c348d4ff",
   135 => x"48c178ff",
   136 => x"f1fd87cb",
   137 => x"058bc187",
   138 => x"c087dbff",
   139 => x"87f1fb48",
   140 => x"5c5b5e0e",
   141 => x"4cd4ff0e",
   142 => x"c687dbfd",
   143 => x"e1c01eea",
   144 => x"49c8c1f0",
   145 => x"c487defb",
   146 => x"02a8c186",
   147 => x"eafe87c8",
   148 => x"c148c087",
   149 => x"dafa87e2",
   150 => x"cf497087",
   151 => x"c699ffff",
   152 => x"c802a9ea",
   153 => x"87d3fe87",
   154 => x"cbc148c0",
   155 => x"7cffc387",
   156 => x"fc4bf1c0",
   157 => x"987087f4",
   158 => x"87ebc002",
   159 => x"ffc01ec0",
   160 => x"49fac1f0",
   161 => x"c487defa",
   162 => x"05987086",
   163 => x"ffc387d9",
   164 => x"c3496c7c",
   165 => x"7c7c7cff",
   166 => x"99c0c17c",
   167 => x"c187c402",
   168 => x"c087d548",
   169 => x"c287d148",
   170 => x"87c405ab",
   171 => x"87c848c0",
   172 => x"fe058bc1",
   173 => x"48c087fd",
   174 => x"1e87e4f9",
   175 => x"dcc21e73",
   176 => x"78c148e0",
   177 => x"d0ff4bc7",
   178 => x"fb78c248",
   179 => x"d0ff87c8",
   180 => x"c078c348",
   181 => x"d0e5c01e",
   182 => x"f949c0c1",
   183 => x"86c487c7",
   184 => x"c105a8c1",
   185 => x"abc24b87",
   186 => x"c087c505",
   187 => x"87f9c048",
   188 => x"ff058bc1",
   189 => x"f7fc87d0",
   190 => x"e4dcc287",
   191 => x"05987058",
   192 => x"1ec187cd",
   193 => x"c1f0ffc0",
   194 => x"d8f849d0",
   195 => x"ff86c487",
   196 => x"ffc348d4",
   197 => x"87e0c478",
   198 => x"58e8dcc2",
   199 => x"c248d0ff",
   200 => x"48d4ff78",
   201 => x"c178ffc3",
   202 => x"87f5f748",
   203 => x"5c5b5e0e",
   204 => x"4a710e5d",
   205 => x"ff4dffc3",
   206 => x"7c754cd4",
   207 => x"c448d0ff",
   208 => x"7c7578c3",
   209 => x"ffc01e72",
   210 => x"49d8c1f0",
   211 => x"c487d6f7",
   212 => x"02987086",
   213 => x"48c087c5",
   214 => x"7587f0c0",
   215 => x"7cfec37c",
   216 => x"d41ec0c8",
   217 => x"dcf54966",
   218 => x"7586c487",
   219 => x"757c757c",
   220 => x"e0dad87c",
   221 => x"6c7c754b",
   222 => x"c5059949",
   223 => x"058bc187",
   224 => x"7c7587f3",
   225 => x"c248d0ff",
   226 => x"f648c178",
   227 => x"ff1e87cf",
   228 => x"d0ff4ad4",
   229 => x"78d1c448",
   230 => x"c17affc3",
   231 => x"87f80589",
   232 => x"731e4f26",
   233 => x"c54b711e",
   234 => x"4adfcdee",
   235 => x"c348d4ff",
   236 => x"486878ff",
   237 => x"02a8fec3",
   238 => x"8ac187c5",
   239 => x"7287ed05",
   240 => x"87c5059a",
   241 => x"eac048c0",
   242 => x"029b7387",
   243 => x"66c887cc",
   244 => x"f449731e",
   245 => x"86c487c5",
   246 => x"66c887c6",
   247 => x"87eefe49",
   248 => x"c348d4ff",
   249 => x"737878ff",
   250 => x"87c5059b",
   251 => x"d048d0ff",
   252 => x"f448c178",
   253 => x"731e87eb",
   254 => x"c04a711e",
   255 => x"48d4ff4b",
   256 => x"ff78ffc3",
   257 => x"c3c448d0",
   258 => x"48d4ff78",
   259 => x"7278ffc3",
   260 => x"f0ffc01e",
   261 => x"f449d1c1",
   262 => x"86c487cb",
   263 => x"cd059870",
   264 => x"1ec0c887",
   265 => x"fd4966cc",
   266 => x"86c487f8",
   267 => x"d0ff4b70",
   268 => x"7378c248",
   269 => x"87e9f348",
   270 => x"5c5b5e0e",
   271 => x"1ec00e5d",
   272 => x"c1f0ffc0",
   273 => x"dcf349c9",
   274 => x"c21ed287",
   275 => x"fd49e8dc",
   276 => x"86c887d0",
   277 => x"84c14cc0",
   278 => x"04acb7d2",
   279 => x"dcc287f8",
   280 => x"49bf97e8",
   281 => x"c199c0c3",
   282 => x"c005a9c0",
   283 => x"dcc287e7",
   284 => x"49bf97ef",
   285 => x"dcc231d0",
   286 => x"4abf97f0",
   287 => x"b17232c8",
   288 => x"97f1dcc2",
   289 => x"71b14abf",
   290 => x"ffffcf4c",
   291 => x"84c19cff",
   292 => x"e7c134ca",
   293 => x"f1dcc287",
   294 => x"c149bf97",
   295 => x"c299c631",
   296 => x"bf97f2dc",
   297 => x"2ab7c74a",
   298 => x"dcc2b172",
   299 => x"4abf97ed",
   300 => x"c29dcf4d",
   301 => x"bf97eedc",
   302 => x"ca9ac34a",
   303 => x"efdcc232",
   304 => x"c24bbf97",
   305 => x"c2b27333",
   306 => x"bf97f0dc",
   307 => x"9bc0c34b",
   308 => x"732bb7c6",
   309 => x"c181c2b2",
   310 => x"70307148",
   311 => x"7548c149",
   312 => x"724d7030",
   313 => x"7184c14c",
   314 => x"b7c0c894",
   315 => x"87cc06ad",
   316 => x"2db734c1",
   317 => x"adb7c0c8",
   318 => x"87f4ff01",
   319 => x"dcf04874",
   320 => x"5b5e0e87",
   321 => x"f80e5d5c",
   322 => x"cee5c286",
   323 => x"c278c048",
   324 => x"c01ec6dd",
   325 => x"87defb49",
   326 => x"987086c4",
   327 => x"c087c505",
   328 => x"87cec948",
   329 => x"7ec14dc0",
   330 => x"bfcbf2c0",
   331 => x"fcddc249",
   332 => x"4bc8714a",
   333 => x"7087f3ec",
   334 => x"87c20598",
   335 => x"f2c07ec0",
   336 => x"c249bfc7",
   337 => x"714ad8de",
   338 => x"ddec4bc8",
   339 => x"05987087",
   340 => x"7ec087c2",
   341 => x"fdc0026e",
   342 => x"cce4c287",
   343 => x"e5c24dbf",
   344 => x"7ebf9fc4",
   345 => x"ead6c548",
   346 => x"87c705a8",
   347 => x"bfcce4c2",
   348 => x"6e87ce4d",
   349 => x"d5e9ca48",
   350 => x"87c502a8",
   351 => x"f1c748c0",
   352 => x"c6ddc287",
   353 => x"f949751e",
   354 => x"86c487ec",
   355 => x"c5059870",
   356 => x"c748c087",
   357 => x"f2c087dc",
   358 => x"c249bfc7",
   359 => x"714ad8de",
   360 => x"c5eb4bc8",
   361 => x"05987087",
   362 => x"e5c287c8",
   363 => x"78c148ce",
   364 => x"f2c087da",
   365 => x"c249bfcb",
   366 => x"714afcdd",
   367 => x"e9ea4bc8",
   368 => x"02987087",
   369 => x"c087c5c0",
   370 => x"87e6c648",
   371 => x"97c4e5c2",
   372 => x"d5c149bf",
   373 => x"cdc005a9",
   374 => x"c5e5c287",
   375 => x"c249bf97",
   376 => x"c002a9ea",
   377 => x"48c087c5",
   378 => x"c287c7c6",
   379 => x"bf97c6dd",
   380 => x"e9c3487e",
   381 => x"cec002a8",
   382 => x"c3486e87",
   383 => x"c002a8eb",
   384 => x"48c087c5",
   385 => x"c287ebc5",
   386 => x"bf97d1dd",
   387 => x"c0059949",
   388 => x"ddc287cc",
   389 => x"49bf97d2",
   390 => x"c002a9c2",
   391 => x"48c087c5",
   392 => x"c287cfc5",
   393 => x"bf97d3dd",
   394 => x"cae5c248",
   395 => x"484c7058",
   396 => x"e5c288c1",
   397 => x"ddc258ce",
   398 => x"49bf97d4",
   399 => x"ddc28175",
   400 => x"4abf97d5",
   401 => x"a17232c8",
   402 => x"dbe9c27e",
   403 => x"c2786e48",
   404 => x"bf97d6dd",
   405 => x"58a6c848",
   406 => x"bfcee5c2",
   407 => x"87d4c202",
   408 => x"bfc7f2c0",
   409 => x"d8dec249",
   410 => x"4bc8714a",
   411 => x"7087fbe7",
   412 => x"c5c00298",
   413 => x"c348c087",
   414 => x"e5c287f8",
   415 => x"c24cbfc6",
   416 => x"c25cefe9",
   417 => x"bf97ebdd",
   418 => x"c231c849",
   419 => x"bf97eadd",
   420 => x"c249a14a",
   421 => x"bf97ecdd",
   422 => x"7232d04a",
   423 => x"ddc249a1",
   424 => x"4abf97ed",
   425 => x"a17232d8",
   426 => x"9166c449",
   427 => x"bfdbe9c2",
   428 => x"e3e9c281",
   429 => x"f3ddc259",
   430 => x"c84abf97",
   431 => x"f2ddc232",
   432 => x"a24bbf97",
   433 => x"f4ddc24a",
   434 => x"d04bbf97",
   435 => x"4aa27333",
   436 => x"97f5ddc2",
   437 => x"9bcf4bbf",
   438 => x"a27333d8",
   439 => x"e7e9c24a",
   440 => x"e3e9c25a",
   441 => x"8ac24abf",
   442 => x"e9c29274",
   443 => x"a17248e7",
   444 => x"87cac178",
   445 => x"97d8ddc2",
   446 => x"31c849bf",
   447 => x"97d7ddc2",
   448 => x"49a14abf",
   449 => x"59d6e5c2",
   450 => x"bfd2e5c2",
   451 => x"c731c549",
   452 => x"29c981ff",
   453 => x"59efe9c2",
   454 => x"97ddddc2",
   455 => x"32c84abf",
   456 => x"97dcddc2",
   457 => x"4aa24bbf",
   458 => x"6e9266c4",
   459 => x"ebe9c282",
   460 => x"e3e9c25a",
   461 => x"c278c048",
   462 => x"7248dfe9",
   463 => x"e9c278a1",
   464 => x"e9c248ef",
   465 => x"c278bfe3",
   466 => x"c248f3e9",
   467 => x"78bfe7e9",
   468 => x"bfcee5c2",
   469 => x"87c9c002",
   470 => x"30c44874",
   471 => x"c9c07e70",
   472 => x"ebe9c287",
   473 => x"30c448bf",
   474 => x"e5c27e70",
   475 => x"786e48d2",
   476 => x"8ef848c1",
   477 => x"4c264d26",
   478 => x"4f264b26",
   479 => x"5c5b5e0e",
   480 => x"4a710e5d",
   481 => x"bfcee5c2",
   482 => x"7287cb02",
   483 => x"722bc74b",
   484 => x"9cffc14c",
   485 => x"4b7287c9",
   486 => x"4c722bc8",
   487 => x"c29cffc3",
   488 => x"83bfdbe9",
   489 => x"bfc3f2c0",
   490 => x"87d902ab",
   491 => x"5bc7f2c0",
   492 => x"1ec6ddc2",
   493 => x"fdf04973",
   494 => x"7086c487",
   495 => x"87c50598",
   496 => x"e6c048c0",
   497 => x"cee5c287",
   498 => x"87d202bf",
   499 => x"91c44974",
   500 => x"81c6ddc2",
   501 => x"ffcf4d69",
   502 => x"9dffffff",
   503 => x"497487cb",
   504 => x"ddc291c2",
   505 => x"699f81c6",
   506 => x"fe48754d",
   507 => x"5e0e87c6",
   508 => x"0e5d5c5b",
   509 => x"c04d711e",
   510 => x"ca49c11e",
   511 => x"86c487ee",
   512 => x"029c4c70",
   513 => x"c287c0c1",
   514 => x"754ad6e5",
   515 => x"87ffe049",
   516 => x"c0029870",
   517 => x"4a7487f1",
   518 => x"4bcb4975",
   519 => x"7087e5e1",
   520 => x"e2c00298",
   521 => x"741ec087",
   522 => x"87c7029c",
   523 => x"c048a6c4",
   524 => x"c487c578",
   525 => x"78c148a6",
   526 => x"c94966c4",
   527 => x"86c487ee",
   528 => x"059c4c70",
   529 => x"7487c0ff",
   530 => x"e7fc2648",
   531 => x"5b5e0e87",
   532 => x"1e0e5d5c",
   533 => x"059b4b71",
   534 => x"48c087c5",
   535 => x"c887e5c1",
   536 => x"7dc04da3",
   537 => x"c70266d4",
   538 => x"9766d487",
   539 => x"87c505bf",
   540 => x"cfc148c0",
   541 => x"4966d487",
   542 => x"7087f3fd",
   543 => x"c1029c4c",
   544 => x"a4dc87c0",
   545 => x"da7d6949",
   546 => x"a3c449a4",
   547 => x"7a699f4a",
   548 => x"bfcee5c2",
   549 => x"d487d202",
   550 => x"699f49a4",
   551 => x"ffffc049",
   552 => x"d0487199",
   553 => x"c27e7030",
   554 => x"6e7ec087",
   555 => x"806a4849",
   556 => x"7bc07a70",
   557 => x"6a49a3cc",
   558 => x"49a3d079",
   559 => x"487479c0",
   560 => x"48c087c2",
   561 => x"87ecfa26",
   562 => x"5c5b5e0e",
   563 => x"4c710e5d",
   564 => x"48c3f2c0",
   565 => x"9c7478ff",
   566 => x"87cac102",
   567 => x"6949a4c8",
   568 => x"87c2c102",
   569 => x"6c4a66d0",
   570 => x"a6d48249",
   571 => x"4d66d05a",
   572 => x"cae5c2b9",
   573 => x"baff4abf",
   574 => x"99719972",
   575 => x"87e4c002",
   576 => x"6b4ba4c4",
   577 => x"87f4f949",
   578 => x"e5c27b70",
   579 => x"6c49bfc6",
   580 => x"757c7181",
   581 => x"cae5c2b9",
   582 => x"baff4abf",
   583 => x"99719972",
   584 => x"87dcff05",
   585 => x"cbf97c75",
   586 => x"1e731e87",
   587 => x"029b4b71",
   588 => x"a3c887c7",
   589 => x"c5056949",
   590 => x"c048c087",
   591 => x"e9c287eb",
   592 => x"c44abfdf",
   593 => x"496949a3",
   594 => x"e5c289c2",
   595 => x"7191bfc6",
   596 => x"e5c24aa2",
   597 => x"6b49bfca",
   598 => x"4aa27199",
   599 => x"721e66c8",
   600 => x"87d2ea49",
   601 => x"497086c4",
   602 => x"87ccf848",
   603 => x"711e731e",
   604 => x"c7029b4b",
   605 => x"49a3c887",
   606 => x"87c50569",
   607 => x"ebc048c0",
   608 => x"dfe9c287",
   609 => x"a3c44abf",
   610 => x"c2496949",
   611 => x"c6e5c289",
   612 => x"a27191bf",
   613 => x"cae5c24a",
   614 => x"996b49bf",
   615 => x"c84aa271",
   616 => x"49721e66",
   617 => x"c487c5e6",
   618 => x"48497086",
   619 => x"0e87c9f7",
   620 => x"5d5c5b5e",
   621 => x"4b711e0e",
   622 => x"c94c66d4",
   623 => x"029b732c",
   624 => x"c887cfc1",
   625 => x"026949a3",
   626 => x"d087c7c1",
   627 => x"66d44da3",
   628 => x"cae5c27d",
   629 => x"b9ff49bf",
   630 => x"7e994a6b",
   631 => x"cd03ac71",
   632 => x"7d7bc087",
   633 => x"c44aa3cc",
   634 => x"796a49a3",
   635 => x"8c7287c2",
   636 => x"dd029c74",
   637 => x"731e4987",
   638 => x"87ccfb49",
   639 => x"66d486c4",
   640 => x"99ffc749",
   641 => x"c287cb02",
   642 => x"731ec6dd",
   643 => x"87d9fc49",
   644 => x"f52686c4",
   645 => x"731e87de",
   646 => x"9b4b711e",
   647 => x"87e4c002",
   648 => x"5bf3e9c2",
   649 => x"8ac24a73",
   650 => x"bfc6e5c2",
   651 => x"e9c29249",
   652 => x"7248bfdf",
   653 => x"f7e9c280",
   654 => x"c4487158",
   655 => x"d6e5c230",
   656 => x"87edc058",
   657 => x"48efe9c2",
   658 => x"bfe3e9c2",
   659 => x"f3e9c278",
   660 => x"e7e9c248",
   661 => x"e5c278bf",
   662 => x"c902bfce",
   663 => x"c6e5c287",
   664 => x"31c449bf",
   665 => x"e9c287c7",
   666 => x"c449bfeb",
   667 => x"d6e5c231",
   668 => x"87c4f459",
   669 => x"5c5b5e0e",
   670 => x"c04a710e",
   671 => x"029a724b",
   672 => x"da87e1c0",
   673 => x"699f49a2",
   674 => x"cee5c24b",
   675 => x"87cf02bf",
   676 => x"9f49a2d4",
   677 => x"c04c4969",
   678 => x"d09cffff",
   679 => x"c087c234",
   680 => x"b349744c",
   681 => x"edfd4973",
   682 => x"87caf387",
   683 => x"5c5b5e0e",
   684 => x"86f40e5d",
   685 => x"7ec04a71",
   686 => x"d8029a72",
   687 => x"c2ddc287",
   688 => x"c278c048",
   689 => x"c248fadc",
   690 => x"78bff3e9",
   691 => x"48fedcc2",
   692 => x"bfefe9c2",
   693 => x"e3e5c278",
   694 => x"c250c048",
   695 => x"49bfd2e5",
   696 => x"bfc2ddc2",
   697 => x"03aa714a",
   698 => x"7287ffc3",
   699 => x"0599cf49",
   700 => x"c287e0c0",
   701 => x"c21ec6dd",
   702 => x"49bffadc",
   703 => x"48fadcc2",
   704 => x"7178a1c1",
   705 => x"c487efe3",
   706 => x"fff1c086",
   707 => x"c6ddc248",
   708 => x"c087cc78",
   709 => x"48bffff1",
   710 => x"c080e0c0",
   711 => x"c258c3f2",
   712 => x"48bfc2dd",
   713 => x"ddc280c1",
   714 => x"7f2758c6",
   715 => x"bf00000c",
   716 => x"9d4dbf97",
   717 => x"87e2c202",
   718 => x"02ade5c3",
   719 => x"c087dbc2",
   720 => x"4bbffff1",
   721 => x"1149a3cb",
   722 => x"05accf4c",
   723 => x"7587d2c1",
   724 => x"c199df49",
   725 => x"c291cd89",
   726 => x"c181d6e5",
   727 => x"51124aa3",
   728 => x"124aa3c3",
   729 => x"4aa3c551",
   730 => x"a3c75112",
   731 => x"c951124a",
   732 => x"51124aa3",
   733 => x"124aa3ce",
   734 => x"4aa3d051",
   735 => x"a3d25112",
   736 => x"d451124a",
   737 => x"51124aa3",
   738 => x"124aa3d6",
   739 => x"4aa3d851",
   740 => x"a3dc5112",
   741 => x"de51124a",
   742 => x"51124aa3",
   743 => x"f9c07ec1",
   744 => x"c8497487",
   745 => x"eac00599",
   746 => x"d0497487",
   747 => x"87d00599",
   748 => x"c00266dc",
   749 => x"497387ca",
   750 => x"700f66dc",
   751 => x"87d30298",
   752 => x"c6c0056e",
   753 => x"d6e5c287",
   754 => x"c050c048",
   755 => x"48bffff1",
   756 => x"c287e7c2",
   757 => x"c048e3e5",
   758 => x"e5c27e50",
   759 => x"c249bfd2",
   760 => x"4abfc2dd",
   761 => x"fc04aa71",
   762 => x"e9c287c1",
   763 => x"c005bff3",
   764 => x"e5c287c8",
   765 => x"c102bfce",
   766 => x"f2c087fe",
   767 => x"78ff48c3",
   768 => x"bffedcc2",
   769 => x"87f4ed49",
   770 => x"ddc24970",
   771 => x"a6c459c2",
   772 => x"fedcc248",
   773 => x"e5c278bf",
   774 => x"c002bfce",
   775 => x"66c487d8",
   776 => x"ffffcf49",
   777 => x"a999f8ff",
   778 => x"87c5c002",
   779 => x"e1c04dc0",
   780 => x"c04dc187",
   781 => x"66c487dc",
   782 => x"f8ffcf49",
   783 => x"c002a999",
   784 => x"a6c887c8",
   785 => x"c078c048",
   786 => x"a6c887c5",
   787 => x"c878c148",
   788 => x"9d754d66",
   789 => x"87e0c005",
   790 => x"c24966c4",
   791 => x"c6e5c289",
   792 => x"c2914abf",
   793 => x"4abfdfe9",
   794 => x"48fadcc2",
   795 => x"c278a172",
   796 => x"c048c2dd",
   797 => x"87e3f978",
   798 => x"8ef448c0",
   799 => x"0087f5eb",
   800 => x"ff000000",
   801 => x"8fffffff",
   802 => x"9800000c",
   803 => x"4600000c",
   804 => x"32335441",
   805 => x"00202020",
   806 => x"31544146",
   807 => x"20202036",
   808 => x"d4ff1e00",
   809 => x"78ffc348",
   810 => x"4f264868",
   811 => x"48d4ff1e",
   812 => x"ff78ffc3",
   813 => x"e1c848d0",
   814 => x"48d4ff78",
   815 => x"e9c278d4",
   816 => x"d4ff48f7",
   817 => x"4f2650bf",
   818 => x"48d0ff1e",
   819 => x"2678e0c0",
   820 => x"ccff1e4f",
   821 => x"99497087",
   822 => x"c087c602",
   823 => x"f105a9fb",
   824 => x"26487187",
   825 => x"5b5e0e4f",
   826 => x"4b710e5c",
   827 => x"f0fe4cc0",
   828 => x"99497087",
   829 => x"87f9c002",
   830 => x"02a9ecc0",
   831 => x"c087f2c0",
   832 => x"c002a9fb",
   833 => x"66cc87eb",
   834 => x"c703acb7",
   835 => x"0266d087",
   836 => x"537187c2",
   837 => x"c2029971",
   838 => x"fe84c187",
   839 => x"497087c3",
   840 => x"87cd0299",
   841 => x"02a9ecc0",
   842 => x"fbc087c7",
   843 => x"d5ff05a9",
   844 => x"0266d087",
   845 => x"97c087c3",
   846 => x"a9ecc07b",
   847 => x"7487c405",
   848 => x"7487c54a",
   849 => x"8a0ac04a",
   850 => x"87c24872",
   851 => x"4c264d26",
   852 => x"4f264b26",
   853 => x"87c9fd1e",
   854 => x"f0c04970",
   855 => x"ca04a9b7",
   856 => x"b7f9c087",
   857 => x"87c301a9",
   858 => x"c189f0c0",
   859 => x"04a9b7c1",
   860 => x"dac187ca",
   861 => x"c301a9b7",
   862 => x"89f7c087",
   863 => x"4f264871",
   864 => x"5c5b5e0e",
   865 => x"ff4a710e",
   866 => x"49724cd4",
   867 => x"7087eac0",
   868 => x"c2029b4b",
   869 => x"ff8bc187",
   870 => x"c5c848d0",
   871 => x"7cd5c178",
   872 => x"31c64973",
   873 => x"97cddbc2",
   874 => x"71484abf",
   875 => x"ff7c70b0",
   876 => x"78c448d0",
   877 => x"d5fe4873",
   878 => x"5b5e0e87",
   879 => x"f80e5d5c",
   880 => x"c04c7186",
   881 => x"87e4fb7e",
   882 => x"f9c04bc0",
   883 => x"49bf97e6",
   884 => x"cf04a9c0",
   885 => x"87f9fb87",
   886 => x"f9c083c1",
   887 => x"49bf97e6",
   888 => x"87f106ab",
   889 => x"97e6f9c0",
   890 => x"87cf02bf",
   891 => x"7087f2fa",
   892 => x"c6029949",
   893 => x"a9ecc087",
   894 => x"c087f105",
   895 => x"87e1fa4b",
   896 => x"dcfa4d70",
   897 => x"58a6c887",
   898 => x"7087d6fa",
   899 => x"c883c14a",
   900 => x"699749a4",
   901 => x"c702ad49",
   902 => x"adffc087",
   903 => x"87e7c005",
   904 => x"9749a4c9",
   905 => x"66c44969",
   906 => x"87c702a9",
   907 => x"a8ffc048",
   908 => x"ca87d405",
   909 => x"699749a4",
   910 => x"c602aa49",
   911 => x"aaffc087",
   912 => x"c187c405",
   913 => x"c087d07e",
   914 => x"c602adec",
   915 => x"adfbc087",
   916 => x"c087c405",
   917 => x"6e7ec14b",
   918 => x"87e1fe02",
   919 => x"7387e9f9",
   920 => x"fb8ef848",
   921 => x"0e0087e6",
   922 => x"5d5c5b5e",
   923 => x"4b711e0e",
   924 => x"ab4d4cc0",
   925 => x"87e8c004",
   926 => x"1ef9f6c0",
   927 => x"c4029d75",
   928 => x"c24ac087",
   929 => x"724ac187",
   930 => x"87e0f049",
   931 => x"7e7086c4",
   932 => x"056e84c1",
   933 => x"4c7387c2",
   934 => x"ac7385c1",
   935 => x"87d8ff06",
   936 => x"2626486e",
   937 => x"264c264d",
   938 => x"0e4f264b",
   939 => x"5d5c5b5e",
   940 => x"4c711e0e",
   941 => x"c291de49",
   942 => x"714dd1ea",
   943 => x"026d9785",
   944 => x"c287ddc1",
   945 => x"4abffce9",
   946 => x"49728274",
   947 => x"7087d8fe",
   948 => x"c0026e7e",
   949 => x"eac287f3",
   950 => x"4a6e4bc4",
   951 => x"c7ff49cb",
   952 => x"4b7487c6",
   953 => x"ddc193cb",
   954 => x"83c483c5",
   955 => x"7be4fcc0",
   956 => x"c2c14974",
   957 => x"7b7587fe",
   958 => x"97d0eac2",
   959 => x"c21e49bf",
   960 => x"c149c4ea",
   961 => x"c487c8de",
   962 => x"c1497486",
   963 => x"c087e5c2",
   964 => x"c4c4c149",
   965 => x"f8e9c287",
   966 => x"c178c048",
   967 => x"87f9dc49",
   968 => x"87fffd26",
   969 => x"64616f4c",
   970 => x"2e676e69",
   971 => x"0e002e2e",
   972 => x"0e5c5b5e",
   973 => x"c24a4b71",
   974 => x"82bffce9",
   975 => x"e6fc4972",
   976 => x"9c4c7087",
   977 => x"4987c402",
   978 => x"c287e9ec",
   979 => x"c048fce9",
   980 => x"dc49c178",
   981 => x"ccfd87c3",
   982 => x"5b5e0e87",
   983 => x"f40e5d5c",
   984 => x"c6ddc286",
   985 => x"c44cc04d",
   986 => x"78c048a6",
   987 => x"bffce9c2",
   988 => x"06a9c049",
   989 => x"c287c1c1",
   990 => x"9848c6dd",
   991 => x"87f8c002",
   992 => x"1ef9f6c0",
   993 => x"c70266c8",
   994 => x"48a6c487",
   995 => x"87c578c0",
   996 => x"c148a6c4",
   997 => x"4966c478",
   998 => x"c487d1ec",
   999 => x"c14d7086",
  1000 => x"4866c484",
  1001 => x"a6c880c1",
  1002 => x"fce9c258",
  1003 => x"03ac49bf",
  1004 => x"9d7587c6",
  1005 => x"87c8ff05",
  1006 => x"9d754cc0",
  1007 => x"87e0c302",
  1008 => x"1ef9f6c0",
  1009 => x"c70266c8",
  1010 => x"48a6cc87",
  1011 => x"87c578c0",
  1012 => x"c148a6cc",
  1013 => x"4966cc78",
  1014 => x"c487d1eb",
  1015 => x"6e7e7086",
  1016 => x"87e9c202",
  1017 => x"81cb496e",
  1018 => x"d0496997",
  1019 => x"d6c10299",
  1020 => x"effcc087",
  1021 => x"cb49744a",
  1022 => x"c5ddc191",
  1023 => x"c8797281",
  1024 => x"51ffc381",
  1025 => x"91de4974",
  1026 => x"4dd1eac2",
  1027 => x"c1c28571",
  1028 => x"a5c17d97",
  1029 => x"51e0c049",
  1030 => x"97d6e5c2",
  1031 => x"87d202bf",
  1032 => x"a5c284c1",
  1033 => x"d6e5c24b",
  1034 => x"ff49db4a",
  1035 => x"c187f9c1",
  1036 => x"a5cd87db",
  1037 => x"c151c049",
  1038 => x"4ba5c284",
  1039 => x"49cb4a6e",
  1040 => x"87e4c1ff",
  1041 => x"c087c6c1",
  1042 => x"744aebfa",
  1043 => x"c191cb49",
  1044 => x"7281c5dd",
  1045 => x"d6e5c279",
  1046 => x"d802bf97",
  1047 => x"de497487",
  1048 => x"c284c191",
  1049 => x"714bd1ea",
  1050 => x"d6e5c283",
  1051 => x"ff49dd4a",
  1052 => x"d887f5c0",
  1053 => x"de4b7487",
  1054 => x"d1eac293",
  1055 => x"49a3cb83",
  1056 => x"84c151c0",
  1057 => x"cb4a6e73",
  1058 => x"dbc0ff49",
  1059 => x"4866c487",
  1060 => x"a6c880c1",
  1061 => x"03acc758",
  1062 => x"6e87c5c0",
  1063 => x"87e0fc05",
  1064 => x"8ef44874",
  1065 => x"1e87fcf7",
  1066 => x"4b711e73",
  1067 => x"c191cb49",
  1068 => x"c881c5dd",
  1069 => x"dbc24aa1",
  1070 => x"501248cd",
  1071 => x"c04aa1c9",
  1072 => x"1248e6f9",
  1073 => x"c281ca50",
  1074 => x"1148d0ea",
  1075 => x"d0eac250",
  1076 => x"1e49bf97",
  1077 => x"d6c149c0",
  1078 => x"e9c287f5",
  1079 => x"78de48f8",
  1080 => x"f4d549c1",
  1081 => x"fef62687",
  1082 => x"4a711e87",
  1083 => x"c191cb49",
  1084 => x"c881c5dd",
  1085 => x"c2481181",
  1086 => x"c258fce9",
  1087 => x"c048fce9",
  1088 => x"d549c178",
  1089 => x"4f2687d3",
  1090 => x"c049c01e",
  1091 => x"2687cafc",
  1092 => x"99711e4f",
  1093 => x"c187d202",
  1094 => x"c048dade",
  1095 => x"c180f750",
  1096 => x"c140e9c3",
  1097 => x"ce78fedc",
  1098 => x"d6dec187",
  1099 => x"f7dcc148",
  1100 => x"c180fc78",
  1101 => x"2678c8c4",
  1102 => x"5b5e0e4f",
  1103 => x"4c710e5c",
  1104 => x"c192cb4a",
  1105 => x"c882c5dd",
  1106 => x"a2c949a2",
  1107 => x"4b6b974b",
  1108 => x"4969971e",
  1109 => x"1282ca1e",
  1110 => x"c5e7c049",
  1111 => x"d349c087",
  1112 => x"497487f7",
  1113 => x"87ccf9c0",
  1114 => x"f8f48ef8",
  1115 => x"1e731e87",
  1116 => x"ff494b71",
  1117 => x"497387c3",
  1118 => x"f487fefe",
  1119 => x"731e87e9",
  1120 => x"c64b711e",
  1121 => x"db024aa3",
  1122 => x"028ac187",
  1123 => x"028a87d6",
  1124 => x"8a87dac1",
  1125 => x"87fcc002",
  1126 => x"e1c0028a",
  1127 => x"cb028a87",
  1128 => x"87dbc187",
  1129 => x"c0fd49c7",
  1130 => x"87dec187",
  1131 => x"bffce9c2",
  1132 => x"87cbc102",
  1133 => x"c288c148",
  1134 => x"c158c0ea",
  1135 => x"eac287c1",
  1136 => x"c002bfc0",
  1137 => x"e9c287f9",
  1138 => x"c148bffc",
  1139 => x"c0eac280",
  1140 => x"87ebc058",
  1141 => x"bffce9c2",
  1142 => x"c289c649",
  1143 => x"c059c0ea",
  1144 => x"da03a9b7",
  1145 => x"fce9c287",
  1146 => x"d278c048",
  1147 => x"c0eac287",
  1148 => x"87cb02bf",
  1149 => x"bffce9c2",
  1150 => x"c280c648",
  1151 => x"c058c0ea",
  1152 => x"87d5d149",
  1153 => x"f6c04973",
  1154 => x"daf287ea",
  1155 => x"5b5e0e87",
  1156 => x"4c710e5c",
  1157 => x"741e66cc",
  1158 => x"c193cb4b",
  1159 => x"c483c5dd",
  1160 => x"496a4aa3",
  1161 => x"87d0fafe",
  1162 => x"7be7c2c1",
  1163 => x"d449a3c8",
  1164 => x"a3c95166",
  1165 => x"5166d849",
  1166 => x"dc49a3ca",
  1167 => x"f1265166",
  1168 => x"5e0e87e3",
  1169 => x"0e5d5c5b",
  1170 => x"d886d0ff",
  1171 => x"a6c459a6",
  1172 => x"c478c048",
  1173 => x"66c4c180",
  1174 => x"c180c478",
  1175 => x"c180c478",
  1176 => x"c0eac278",
  1177 => x"c278c148",
  1178 => x"48bff8e9",
  1179 => x"cb05a8de",
  1180 => x"87e5f387",
  1181 => x"a6c84970",
  1182 => x"87e6ce59",
  1183 => x"e987ede8",
  1184 => x"dce887cf",
  1185 => x"c04c7087",
  1186 => x"c102acfb",
  1187 => x"66d487d0",
  1188 => x"87c2c105",
  1189 => x"c11e1ec0",
  1190 => x"f8dec11e",
  1191 => x"fd49c01e",
  1192 => x"d0c187eb",
  1193 => x"82c44a66",
  1194 => x"81c7496a",
  1195 => x"1ec15174",
  1196 => x"496a1ed8",
  1197 => x"ece881c8",
  1198 => x"c186d887",
  1199 => x"c04866c4",
  1200 => x"87c701a8",
  1201 => x"c148a6c4",
  1202 => x"c187ce78",
  1203 => x"c14866c4",
  1204 => x"58a6cc88",
  1205 => x"f8e787c3",
  1206 => x"48a6cc87",
  1207 => x"9c7478c2",
  1208 => x"87facc02",
  1209 => x"c14866c4",
  1210 => x"03a866c8",
  1211 => x"d887efcc",
  1212 => x"78c048a6",
  1213 => x"78c080c4",
  1214 => x"7087e6e6",
  1215 => x"acd0c14c",
  1216 => x"87d7c205",
  1217 => x"e97e66dc",
  1218 => x"497087ca",
  1219 => x"59a6e0c0",
  1220 => x"7087cee6",
  1221 => x"acecc04c",
  1222 => x"87eac105",
  1223 => x"cb4966c4",
  1224 => x"66c0c191",
  1225 => x"4aa1c481",
  1226 => x"a1c84d6a",
  1227 => x"5266dc4a",
  1228 => x"79e9c3c1",
  1229 => x"7087eae5",
  1230 => x"d8029c4c",
  1231 => x"acfbc087",
  1232 => x"7487d202",
  1233 => x"87d9e555",
  1234 => x"029c4c70",
  1235 => x"fbc087c7",
  1236 => x"eeff05ac",
  1237 => x"55e0c087",
  1238 => x"c055c1c2",
  1239 => x"66d47d97",
  1240 => x"05a96e49",
  1241 => x"66c487db",
  1242 => x"a866c848",
  1243 => x"c487ca04",
  1244 => x"80c14866",
  1245 => x"c858a6c8",
  1246 => x"4866c887",
  1247 => x"a6cc88c1",
  1248 => x"87dde458",
  1249 => x"d0c14c70",
  1250 => x"87c805ac",
  1251 => x"c14866d0",
  1252 => x"58a6d480",
  1253 => x"02acd0c1",
  1254 => x"c087e9fd",
  1255 => x"d448a6e0",
  1256 => x"66dc7866",
  1257 => x"66e0c048",
  1258 => x"c3c905a8",
  1259 => x"a6e4c087",
  1260 => x"7e78c048",
  1261 => x"fbc04874",
  1262 => x"a6ecc088",
  1263 => x"02987058",
  1264 => x"4887c8c8",
  1265 => x"ecc088cb",
  1266 => x"987058a6",
  1267 => x"87d0c102",
  1268 => x"c088c948",
  1269 => x"7058a6ec",
  1270 => x"d6c30298",
  1271 => x"88c44887",
  1272 => x"58a6ecc0",
  1273 => x"d0029870",
  1274 => x"88c14887",
  1275 => x"58a6ecc0",
  1276 => x"c2029870",
  1277 => x"ccc787fd",
  1278 => x"48a6d887",
  1279 => x"e278f0c0",
  1280 => x"4c7087df",
  1281 => x"02acecc0",
  1282 => x"dc87c3c0",
  1283 => x"ecc05ca6",
  1284 => x"87cc02ac",
  1285 => x"7087cae2",
  1286 => x"acecc04c",
  1287 => x"87f4ff05",
  1288 => x"02acecc0",
  1289 => x"e187c3c0",
  1290 => x"66d887f7",
  1291 => x"4966d41e",
  1292 => x"4966d41e",
  1293 => x"f8dec11e",
  1294 => x"4966d41e",
  1295 => x"c087cef7",
  1296 => x"dc1eca1e",
  1297 => x"91cb4966",
  1298 => x"8166d8c1",
  1299 => x"c448a6d8",
  1300 => x"66d878a1",
  1301 => x"cce249bf",
  1302 => x"c086d887",
  1303 => x"c106a8b7",
  1304 => x"1ec187c4",
  1305 => x"66c81ede",
  1306 => x"f8e149bf",
  1307 => x"7086c887",
  1308 => x"08c04849",
  1309 => x"58a6dc88",
  1310 => x"06a8b7c0",
  1311 => x"d887e7c0",
  1312 => x"b7dd4866",
  1313 => x"87de03a8",
  1314 => x"d849bf6e",
  1315 => x"e0c08166",
  1316 => x"4966d851",
  1317 => x"bf6e81c1",
  1318 => x"51c1c281",
  1319 => x"c24966d8",
  1320 => x"81bf6e81",
  1321 => x"66cc51c0",
  1322 => x"d080c148",
  1323 => x"7ec158a6",
  1324 => x"e287d8c4",
  1325 => x"a6dc87de",
  1326 => x"87d8e258",
  1327 => x"58a6ecc0",
  1328 => x"05a8ecc0",
  1329 => x"c087cac0",
  1330 => x"d848a6e8",
  1331 => x"c4c07866",
  1332 => x"ccdfff87",
  1333 => x"4966c487",
  1334 => x"c0c191cb",
  1335 => x"80714866",
  1336 => x"4a6e7e70",
  1337 => x"496e82c8",
  1338 => x"66d881ca",
  1339 => x"66e8c051",
  1340 => x"d881c149",
  1341 => x"48c18966",
  1342 => x"49703071",
  1343 => x"977189c1",
  1344 => x"ededc27a",
  1345 => x"66d849bf",
  1346 => x"4a6a9729",
  1347 => x"c0987148",
  1348 => x"6e58a6f0",
  1349 => x"6981c449",
  1350 => x"66e0c04d",
  1351 => x"a866dc48",
  1352 => x"87c8c002",
  1353 => x"c048a6d8",
  1354 => x"87c5c078",
  1355 => x"c148a6d8",
  1356 => x"1e66d878",
  1357 => x"751ee0c0",
  1358 => x"e8deff49",
  1359 => x"7086c887",
  1360 => x"acb7c04c",
  1361 => x"87d4c106",
  1362 => x"e0c08574",
  1363 => x"75897449",
  1364 => x"d6d9c14b",
  1365 => x"edfe714a",
  1366 => x"85c287ce",
  1367 => x"4866e4c0",
  1368 => x"e8c080c1",
  1369 => x"ecc058a6",
  1370 => x"81c14966",
  1371 => x"c002a970",
  1372 => x"a6d887c8",
  1373 => x"c078c048",
  1374 => x"a6d887c5",
  1375 => x"d878c148",
  1376 => x"a4c21e66",
  1377 => x"48e0c049",
  1378 => x"49708871",
  1379 => x"ff49751e",
  1380 => x"c887d2dd",
  1381 => x"a8b7c086",
  1382 => x"87c0ff01",
  1383 => x"0266e4c0",
  1384 => x"6e87d1c0",
  1385 => x"c081c949",
  1386 => x"6e5166e4",
  1387 => x"f9c4c148",
  1388 => x"87ccc078",
  1389 => x"81c9496e",
  1390 => x"486e51c2",
  1391 => x"78edc5c1",
  1392 => x"c6c07ec1",
  1393 => x"c8dcff87",
  1394 => x"6e4c7087",
  1395 => x"87f5c002",
  1396 => x"c84866c4",
  1397 => x"c004a866",
  1398 => x"66c487cb",
  1399 => x"c880c148",
  1400 => x"e0c058a6",
  1401 => x"4866c887",
  1402 => x"a6cc88c1",
  1403 => x"87d5c058",
  1404 => x"05acc6c1",
  1405 => x"cc87c8c0",
  1406 => x"80c14866",
  1407 => x"ff58a6d0",
  1408 => x"7087cedb",
  1409 => x"4866d04c",
  1410 => x"a6d480c1",
  1411 => x"029c7458",
  1412 => x"c487cbc0",
  1413 => x"c8c14866",
  1414 => x"f304a866",
  1415 => x"daff87d1",
  1416 => x"66c487e6",
  1417 => x"03a8c748",
  1418 => x"c287e5c0",
  1419 => x"c048c0ea",
  1420 => x"4966c478",
  1421 => x"c0c191cb",
  1422 => x"a1c48166",
  1423 => x"c04a6a4a",
  1424 => x"66c47952",
  1425 => x"c880c148",
  1426 => x"a8c758a6",
  1427 => x"87dbff04",
  1428 => x"e18ed0ff",
  1429 => x"203a87cd",
  1430 => x"1e731e00",
  1431 => x"029b4b71",
  1432 => x"e9c287c6",
  1433 => x"78c048fc",
  1434 => x"e9c21ec7",
  1435 => x"1e49bffc",
  1436 => x"1ec5ddc1",
  1437 => x"bff8e9c2",
  1438 => x"87c6ef49",
  1439 => x"e9c286cc",
  1440 => x"ea49bff8",
  1441 => x"9b7387cb",
  1442 => x"c187c802",
  1443 => x"c049c5dd",
  1444 => x"e087f3e5",
  1445 => x"c21e87d1",
  1446 => x"c048cddb",
  1447 => x"e8dec150",
  1448 => x"fbc049bf",
  1449 => x"48c087fc",
  1450 => x"c71e4f26",
  1451 => x"49c187e9",
  1452 => x"fe87e6fe",
  1453 => x"7087c4f0",
  1454 => x"87cd0298",
  1455 => x"87c1f9fe",
  1456 => x"c4029870",
  1457 => x"c24ac187",
  1458 => x"724ac087",
  1459 => x"87ce059a",
  1460 => x"dbc11ec0",
  1461 => x"f1c049fe",
  1462 => x"86c487f0",
  1463 => x"c0c187fe",
  1464 => x"1ec087d5",
  1465 => x"49c9dcc1",
  1466 => x"87def1c0",
  1467 => x"e5fe1ec0",
  1468 => x"c0497087",
  1469 => x"c387d3f1",
  1470 => x"8ef887dc",
  1471 => x"44534f26",
  1472 => x"69616620",
  1473 => x"2e64656c",
  1474 => x"6f6f4200",
  1475 => x"676e6974",
  1476 => x"002e2e2e",
  1477 => x"c9e8c01e",
  1478 => x"f4f4c087",
  1479 => x"2687f687",
  1480 => x"e9c21e4f",
  1481 => x"78c048fc",
  1482 => x"48f8e9c2",
  1483 => x"f9fd78c0",
  1484 => x"c087e187",
  1485 => x"804f2648",
  1486 => x"69784520",
  1487 => x"20800074",
  1488 => x"6b636142",
  1489 => x"0010e900",
  1490 => x"002a9100",
  1491 => x"00000000",
  1492 => x"000010e9",
  1493 => x"00002aaf",
  1494 => x"e9000000",
  1495 => x"cd000010",
  1496 => x"0000002a",
  1497 => x"10e90000",
  1498 => x"2aeb0000",
  1499 => x"00000000",
  1500 => x"0010e900",
  1501 => x"002b0900",
  1502 => x"00000000",
  1503 => x"000010e9",
  1504 => x"00002b27",
  1505 => x"e9000000",
  1506 => x"45000010",
  1507 => x"0000002b",
  1508 => x"10e90000",
  1509 => x"00000000",
  1510 => x"00000000",
  1511 => x"00117e00",
  1512 => x"00000000",
  1513 => x"00000000",
  1514 => x"000017ac",
  1515 => x"544f4f42",
  1516 => x"20202020",
  1517 => x"004d4f52",
  1518 => x"64616f4c",
  1519 => x"002e2a20",
  1520 => x"48f0fe1e",
  1521 => x"09cd78c0",
  1522 => x"4f260979",
  1523 => x"f0fe1e1e",
  1524 => x"26487ebf",
  1525 => x"fe1e4f26",
  1526 => x"78c148f0",
  1527 => x"fe1e4f26",
  1528 => x"78c048f0",
  1529 => x"711e4f26",
  1530 => x"5252c04a",
  1531 => x"5e0e4f26",
  1532 => x"0e5d5c5b",
  1533 => x"4d7186f4",
  1534 => x"c17e6d97",
  1535 => x"6c974ca5",
  1536 => x"58a6c848",
  1537 => x"66c4486e",
  1538 => x"87c505a8",
  1539 => x"e6c048ff",
  1540 => x"87caff87",
  1541 => x"9749a5c2",
  1542 => x"a3714b6c",
  1543 => x"4b6b974b",
  1544 => x"6e7e6c97",
  1545 => x"c880c148",
  1546 => x"98c758a6",
  1547 => x"7058a6cc",
  1548 => x"e1fe7c97",
  1549 => x"f4487387",
  1550 => x"264d268e",
  1551 => x"264b264c",
  1552 => x"5b5e0e4f",
  1553 => x"86f40e5c",
  1554 => x"66d84c71",
  1555 => x"9affc34a",
  1556 => x"974ba4c2",
  1557 => x"a173496c",
  1558 => x"97517249",
  1559 => x"486e7e6c",
  1560 => x"a6c880c1",
  1561 => x"cc98c758",
  1562 => x"547058a6",
  1563 => x"caff8ef4",
  1564 => x"fd1e1e87",
  1565 => x"bfe087e8",
  1566 => x"e0c0494a",
  1567 => x"cb0299c0",
  1568 => x"c21e7287",
  1569 => x"fe49e3ed",
  1570 => x"86c487f7",
  1571 => x"7087fdfc",
  1572 => x"87c2fd7e",
  1573 => x"1e4f2626",
  1574 => x"49e3edc2",
  1575 => x"c187c7fd",
  1576 => x"fc49f1e1",
  1577 => x"d9c587da",
  1578 => x"0e4f2687",
  1579 => x"5d5c5b5e",
  1580 => x"c2eec20e",
  1581 => x"e3c14abf",
  1582 => x"4c49bfff",
  1583 => x"4d71bc72",
  1584 => x"c087dbfc",
  1585 => x"d049744b",
  1586 => x"87d50299",
  1587 => x"99d04975",
  1588 => x"1ec01e71",
  1589 => x"4ad1eac1",
  1590 => x"49128273",
  1591 => x"c887e4c0",
  1592 => x"2d2cc186",
  1593 => x"04abc883",
  1594 => x"fb87daff",
  1595 => x"e3c187e8",
  1596 => x"eec248ff",
  1597 => x"2678bfc2",
  1598 => x"264c264d",
  1599 => x"004f264b",
  1600 => x"1e000000",
  1601 => x"c848d0ff",
  1602 => x"d4ff78e1",
  1603 => x"c478c548",
  1604 => x"87c30266",
  1605 => x"c878e0c3",
  1606 => x"87c60266",
  1607 => x"c348d4ff",
  1608 => x"d4ff78f0",
  1609 => x"ff787148",
  1610 => x"e1c848d0",
  1611 => x"78e0c078",
  1612 => x"5e0e4f26",
  1613 => x"710e5c5b",
  1614 => x"e3edc24c",
  1615 => x"87eefa49",
  1616 => x"b7c04a70",
  1617 => x"e3c204aa",
  1618 => x"aae0c387",
  1619 => x"c187c905",
  1620 => x"c148f5e7",
  1621 => x"87d4c278",
  1622 => x"05aaf0c3",
  1623 => x"e7c187c9",
  1624 => x"78c148f1",
  1625 => x"c187f5c1",
  1626 => x"02bff5e7",
  1627 => x"4b7287c7",
  1628 => x"c2b3c0c2",
  1629 => x"744b7287",
  1630 => x"87d1059c",
  1631 => x"bff1e7c1",
  1632 => x"f5e7c11e",
  1633 => x"49721ebf",
  1634 => x"c887f8fd",
  1635 => x"f1e7c186",
  1636 => x"e0c002bf",
  1637 => x"c4497387",
  1638 => x"c19129b7",
  1639 => x"7381d1e9",
  1640 => x"c29acf4a",
  1641 => x"7248c192",
  1642 => x"ff4a7030",
  1643 => x"694872ba",
  1644 => x"db797098",
  1645 => x"c4497387",
  1646 => x"c19129b7",
  1647 => x"7381d1e9",
  1648 => x"c29acf4a",
  1649 => x"7248c392",
  1650 => x"484a7030",
  1651 => x"7970b069",
  1652 => x"48f5e7c1",
  1653 => x"e7c178c0",
  1654 => x"78c048f1",
  1655 => x"49e3edc2",
  1656 => x"7087cbf8",
  1657 => x"aab7c04a",
  1658 => x"87ddfd03",
  1659 => x"c8fc48c0",
  1660 => x"00000087",
  1661 => x"00000000",
  1662 => x"4a711e00",
  1663 => x"87f2fc49",
  1664 => x"c01e4f26",
  1665 => x"c449724a",
  1666 => x"d1e9c191",
  1667 => x"c179c081",
  1668 => x"aab7d082",
  1669 => x"2687ee04",
  1670 => x"5b5e0e4f",
  1671 => x"710e5d5c",
  1672 => x"87faf64d",
  1673 => x"b7c44a75",
  1674 => x"e9c1922a",
  1675 => x"4c7582d1",
  1676 => x"94c29ccf",
  1677 => x"744b496a",
  1678 => x"c29bc32b",
  1679 => x"70307448",
  1680 => x"74bcff4c",
  1681 => x"70987148",
  1682 => x"87caf67a",
  1683 => x"e6fa4873",
  1684 => x"00000087",
  1685 => x"00000000",
  1686 => x"00000000",
  1687 => x"00000000",
  1688 => x"00000000",
  1689 => x"00000000",
  1690 => x"00000000",
  1691 => x"00000000",
  1692 => x"00000000",
  1693 => x"00000000",
  1694 => x"00000000",
  1695 => x"00000000",
  1696 => x"00000000",
  1697 => x"00000000",
  1698 => x"00000000",
  1699 => x"00000000",
  1700 => x"261e1600",
  1701 => x"3d362e25",
  1702 => x"d0ff1e3e",
  1703 => x"78e1c848",
  1704 => x"d4ff4871",
  1705 => x"4f267808",
  1706 => x"48d0ff1e",
  1707 => x"7178e1c8",
  1708 => x"08d4ff48",
  1709 => x"4866c478",
  1710 => x"7808d4ff",
  1711 => x"711e4f26",
  1712 => x"4966c44a",
  1713 => x"ff49721e",
  1714 => x"d0ff87de",
  1715 => x"78e0c048",
  1716 => x"1e4f2626",
  1717 => x"66c44a71",
  1718 => x"a2e0c11e",
  1719 => x"87c8ff49",
  1720 => x"c84966c8",
  1721 => x"d4ff29b7",
  1722 => x"ff787148",
  1723 => x"e0c048d0",
  1724 => x"4f262678",
  1725 => x"4ad4ff1e",
  1726 => x"ff7affc3",
  1727 => x"e1c848d0",
  1728 => x"c27ade78",
  1729 => x"7abfeded",
  1730 => x"28c84849",
  1731 => x"48717a70",
  1732 => x"7a7028d0",
  1733 => x"28d84871",
  1734 => x"d0ff7a70",
  1735 => x"78e0c048",
  1736 => x"5e0e4f26",
  1737 => x"0e5d5c5b",
  1738 => x"edc24c71",
  1739 => x"4b4dbfed",
  1740 => x"66d02b74",
  1741 => x"d483c19b",
  1742 => x"c204ab66",
  1743 => x"744bc087",
  1744 => x"4966d04a",
  1745 => x"b9ff3172",
  1746 => x"48739975",
  1747 => x"4a703072",
  1748 => x"c2b07148",
  1749 => x"fe58f1ed",
  1750 => x"4d2687da",
  1751 => x"4b264c26",
  1752 => x"ff1e4f26",
  1753 => x"c9c848d0",
  1754 => x"ff487178",
  1755 => x"267808d4",
  1756 => x"4a711e4f",
  1757 => x"ff87eb49",
  1758 => x"78c848d0",
  1759 => x"731e4f26",
  1760 => x"c24b711e",
  1761 => x"02bffded",
  1762 => x"ebc287c3",
  1763 => x"48d0ff87",
  1764 => x"7378c9c8",
  1765 => x"b1e0c049",
  1766 => x"7148d4ff",
  1767 => x"f1edc278",
  1768 => x"c878c048",
  1769 => x"87c50266",
  1770 => x"c249ffc3",
  1771 => x"c249c087",
  1772 => x"cc59f9ed",
  1773 => x"87c60266",
  1774 => x"4ad5d5c5",
  1775 => x"ffcf87c4",
  1776 => x"edc24aff",
  1777 => x"edc25afd",
  1778 => x"78c148fd",
  1779 => x"4d2687c4",
  1780 => x"4b264c26",
  1781 => x"5e0e4f26",
  1782 => x"0e5d5c5b",
  1783 => x"edc24a71",
  1784 => x"724cbff9",
  1785 => x"87cb029a",
  1786 => x"c191c849",
  1787 => x"714bf4ed",
  1788 => x"c187c483",
  1789 => x"c04bf4f1",
  1790 => x"7449134d",
  1791 => x"f5edc299",
  1792 => x"d4ffb9bf",
  1793 => x"c1787148",
  1794 => x"c8852cb7",
  1795 => x"e804adb7",
  1796 => x"f1edc287",
  1797 => x"80c848bf",
  1798 => x"58f5edc2",
  1799 => x"1e87effe",
  1800 => x"4b711e73",
  1801 => x"029a4a13",
  1802 => x"497287cb",
  1803 => x"1387e7fe",
  1804 => x"f5059a4a",
  1805 => x"87dafe87",
  1806 => x"f1edc21e",
  1807 => x"edc249bf",
  1808 => x"a1c148f1",
  1809 => x"b7c0c478",
  1810 => x"87db03a9",
  1811 => x"c248d4ff",
  1812 => x"78bff5ed",
  1813 => x"bff1edc2",
  1814 => x"f1edc249",
  1815 => x"78a1c148",
  1816 => x"a9b7c0c4",
  1817 => x"ff87e504",
  1818 => x"78c848d0",
  1819 => x"48fdedc2",
  1820 => x"4f2678c0",
  1821 => x"00000000",
  1822 => x"00000000",
  1823 => x"5f000000",
  1824 => x"0000005f",
  1825 => x"00030300",
  1826 => x"00000303",
  1827 => x"147f7f14",
  1828 => x"00147f7f",
  1829 => x"6b2e2400",
  1830 => x"00123a6b",
  1831 => x"18366a4c",
  1832 => x"0032566c",
  1833 => x"594f7e30",
  1834 => x"40683a77",
  1835 => x"07040000",
  1836 => x"00000003",
  1837 => x"3e1c0000",
  1838 => x"00004163",
  1839 => x"63410000",
  1840 => x"00001c3e",
  1841 => x"1c3e2a08",
  1842 => x"082a3e1c",
  1843 => x"3e080800",
  1844 => x"0008083e",
  1845 => x"e0800000",
  1846 => x"00000060",
  1847 => x"08080800",
  1848 => x"00080808",
  1849 => x"60000000",
  1850 => x"00000060",
  1851 => x"18306040",
  1852 => x"0103060c",
  1853 => x"597f3e00",
  1854 => x"003e7f4d",
  1855 => x"7f060400",
  1856 => x"0000007f",
  1857 => x"71634200",
  1858 => x"00464f59",
  1859 => x"49632200",
  1860 => x"00367f49",
  1861 => x"13161c18",
  1862 => x"00107f7f",
  1863 => x"45672700",
  1864 => x"00397d45",
  1865 => x"4b7e3c00",
  1866 => x"00307949",
  1867 => x"71010100",
  1868 => x"00070f79",
  1869 => x"497f3600",
  1870 => x"00367f49",
  1871 => x"494f0600",
  1872 => x"001e3f69",
  1873 => x"66000000",
  1874 => x"00000066",
  1875 => x"e6800000",
  1876 => x"00000066",
  1877 => x"14080800",
  1878 => x"00222214",
  1879 => x"14141400",
  1880 => x"00141414",
  1881 => x"14222200",
  1882 => x"00080814",
  1883 => x"51030200",
  1884 => x"00060f59",
  1885 => x"5d417f3e",
  1886 => x"001e1f55",
  1887 => x"097f7e00",
  1888 => x"007e7f09",
  1889 => x"497f7f00",
  1890 => x"00367f49",
  1891 => x"633e1c00",
  1892 => x"00414141",
  1893 => x"417f7f00",
  1894 => x"001c3e63",
  1895 => x"497f7f00",
  1896 => x"00414149",
  1897 => x"097f7f00",
  1898 => x"00010109",
  1899 => x"417f3e00",
  1900 => x"007a7b49",
  1901 => x"087f7f00",
  1902 => x"007f7f08",
  1903 => x"7f410000",
  1904 => x"0000417f",
  1905 => x"40602000",
  1906 => x"003f7f40",
  1907 => x"1c087f7f",
  1908 => x"00416336",
  1909 => x"407f7f00",
  1910 => x"00404040",
  1911 => x"0c067f7f",
  1912 => x"007f7f06",
  1913 => x"0c067f7f",
  1914 => x"007f7f18",
  1915 => x"417f3e00",
  1916 => x"003e7f41",
  1917 => x"097f7f00",
  1918 => x"00060f09",
  1919 => x"61417f3e",
  1920 => x"00407e7f",
  1921 => x"097f7f00",
  1922 => x"00667f19",
  1923 => x"4d6f2600",
  1924 => x"00327b59",
  1925 => x"7f010100",
  1926 => x"0001017f",
  1927 => x"407f3f00",
  1928 => x"003f7f40",
  1929 => x"703f0f00",
  1930 => x"000f3f70",
  1931 => x"18307f7f",
  1932 => x"007f7f30",
  1933 => x"1c366341",
  1934 => x"4163361c",
  1935 => x"7c060301",
  1936 => x"0103067c",
  1937 => x"4d597161",
  1938 => x"00414347",
  1939 => x"7f7f0000",
  1940 => x"00004141",
  1941 => x"0c060301",
  1942 => x"40603018",
  1943 => x"41410000",
  1944 => x"00007f7f",
  1945 => x"03060c08",
  1946 => x"00080c06",
  1947 => x"80808080",
  1948 => x"00808080",
  1949 => x"03000000",
  1950 => x"00000407",
  1951 => x"54742000",
  1952 => x"00787c54",
  1953 => x"447f7f00",
  1954 => x"00387c44",
  1955 => x"447c3800",
  1956 => x"00004444",
  1957 => x"447c3800",
  1958 => x"007f7f44",
  1959 => x"547c3800",
  1960 => x"00185c54",
  1961 => x"7f7e0400",
  1962 => x"00000505",
  1963 => x"a4bc1800",
  1964 => x"007cfca4",
  1965 => x"047f7f00",
  1966 => x"00787c04",
  1967 => x"3d000000",
  1968 => x"0000407d",
  1969 => x"80808000",
  1970 => x"00007dfd",
  1971 => x"107f7f00",
  1972 => x"00446c38",
  1973 => x"3f000000",
  1974 => x"0000407f",
  1975 => x"180c7c7c",
  1976 => x"00787c0c",
  1977 => x"047c7c00",
  1978 => x"00787c04",
  1979 => x"447c3800",
  1980 => x"00387c44",
  1981 => x"24fcfc00",
  1982 => x"00183c24",
  1983 => x"243c1800",
  1984 => x"00fcfc24",
  1985 => x"047c7c00",
  1986 => x"00080c04",
  1987 => x"545c4800",
  1988 => x"00207454",
  1989 => x"7f3f0400",
  1990 => x"00004444",
  1991 => x"407c3c00",
  1992 => x"007c7c40",
  1993 => x"603c1c00",
  1994 => x"001c3c60",
  1995 => x"30607c3c",
  1996 => x"003c7c60",
  1997 => x"10386c44",
  1998 => x"00446c38",
  1999 => x"e0bc1c00",
  2000 => x"001c3c60",
  2001 => x"74644400",
  2002 => x"00444c5c",
  2003 => x"3e080800",
  2004 => x"00414177",
  2005 => x"7f000000",
  2006 => x"0000007f",
  2007 => x"77414100",
  2008 => x"0008083e",
  2009 => x"03010102",
  2010 => x"00010202",
  2011 => x"7f7f7f7f",
  2012 => x"007f7f7f",
  2013 => x"1c1c0808",
  2014 => x"7f7f3e3e",
  2015 => x"3e3e7f7f",
  2016 => x"08081c1c",
  2017 => x"7c181000",
  2018 => x"0010187c",
  2019 => x"7c301000",
  2020 => x"0010307c",
  2021 => x"60603010",
  2022 => x"00061e78",
  2023 => x"183c6642",
  2024 => x"0042663c",
  2025 => x"c26a3878",
  2026 => x"00386cc6",
  2027 => x"60000060",
  2028 => x"00600000",
  2029 => x"5c5b5e0e",
  2030 => x"711e0e5d",
  2031 => x"ceeec24c",
  2032 => x"4bc04dbf",
  2033 => x"ab741ec0",
  2034 => x"c487c702",
  2035 => x"78c048a6",
  2036 => x"a6c487c5",
  2037 => x"c478c148",
  2038 => x"49731e66",
  2039 => x"c887dfee",
  2040 => x"49e0c086",
  2041 => x"c487efef",
  2042 => x"496a4aa5",
  2043 => x"f187f0f0",
  2044 => x"85cb87c6",
  2045 => x"b7c883c1",
  2046 => x"c7ff04ab",
  2047 => x"4d262687",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
