
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"d4",x"ef",x"c2",x"87"),
    12 => (x"86",x"c0",x"c6",x"4e"),
    13 => (x"49",x"d4",x"ef",x"c2"),
    14 => (x"48",x"e0",x"dc",x"c2"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"d6",x"db"),
    19 => (x"1e",x"87",x"fc",x"98"),
    20 => (x"1e",x"73",x"1e",x"72"),
    21 => (x"02",x"11",x"48",x"12"),
    22 => (x"c3",x"4b",x"87",x"ca"),
    23 => (x"73",x"9b",x"98",x"df"),
    24 => (x"87",x"f0",x"02",x"88"),
    25 => (x"4a",x"26",x"4b",x"26"),
    26 => (x"73",x"1e",x"4f",x"26"),
    27 => (x"c1",x"1e",x"72",x"1e"),
    28 => (x"87",x"ca",x"04",x"8b"),
    29 => (x"02",x"11",x"48",x"12"),
    30 => (x"02",x"88",x"87",x"c4"),
    31 => (x"4a",x"26",x"87",x"f1"),
    32 => (x"4f",x"26",x"4b",x"26"),
    33 => (x"73",x"1e",x"74",x"1e"),
    34 => (x"c1",x"1e",x"72",x"1e"),
    35 => (x"87",x"d0",x"04",x"8b"),
    36 => (x"02",x"11",x"48",x"12"),
    37 => (x"c3",x"4c",x"87",x"ca"),
    38 => (x"74",x"9c",x"98",x"df"),
    39 => (x"87",x"eb",x"02",x"88"),
    40 => (x"4b",x"26",x"4a",x"26"),
    41 => (x"4f",x"26",x"4c",x"26"),
    42 => (x"81",x"48",x"73",x"1e"),
    43 => (x"c5",x"02",x"a9",x"73"),
    44 => (x"05",x"53",x"12",x"87"),
    45 => (x"4f",x"26",x"87",x"f6"),
    46 => (x"4a",x"66",x"c4",x"1e"),
    47 => (x"51",x"12",x"48",x"71"),
    48 => (x"26",x"87",x"fb",x"05"),
    49 => (x"48",x"11",x"1e",x"4f"),
    50 => (x"78",x"08",x"d4",x"ff"),
    51 => (x"c1",x"48",x"66",x"c4"),
    52 => (x"58",x"a6",x"c8",x"88"),
    53 => (x"ed",x"05",x"98",x"70"),
    54 => (x"1e",x"4f",x"26",x"87"),
    55 => (x"c3",x"48",x"d4",x"ff"),
    56 => (x"51",x"68",x"78",x"ff"),
    57 => (x"c1",x"48",x"66",x"c4"),
    58 => (x"58",x"a6",x"c8",x"88"),
    59 => (x"eb",x"05",x"98",x"70"),
    60 => (x"1e",x"4f",x"26",x"87"),
    61 => (x"d4",x"ff",x"1e",x"73"),
    62 => (x"7b",x"ff",x"c3",x"4b"),
    63 => (x"ff",x"c3",x"4a",x"6b"),
    64 => (x"c8",x"49",x"6b",x"7b"),
    65 => (x"c3",x"b1",x"72",x"32"),
    66 => (x"4a",x"6b",x"7b",x"ff"),
    67 => (x"b2",x"71",x"31",x"c8"),
    68 => (x"6b",x"7b",x"ff",x"c3"),
    69 => (x"72",x"32",x"c8",x"49"),
    70 => (x"c4",x"48",x"71",x"b1"),
    71 => (x"26",x"4d",x"26",x"87"),
    72 => (x"26",x"4b",x"26",x"4c"),
    73 => (x"5b",x"5e",x"0e",x"4f"),
    74 => (x"71",x"0e",x"5d",x"5c"),
    75 => (x"4c",x"d4",x"ff",x"4a"),
    76 => (x"ff",x"c3",x"49",x"72"),
    77 => (x"c2",x"7c",x"71",x"99"),
    78 => (x"05",x"bf",x"e0",x"dc"),
    79 => (x"66",x"d0",x"87",x"c8"),
    80 => (x"d4",x"30",x"c9",x"48"),
    81 => (x"66",x"d0",x"58",x"a6"),
    82 => (x"c3",x"29",x"d8",x"49"),
    83 => (x"7c",x"71",x"99",x"ff"),
    84 => (x"d0",x"49",x"66",x"d0"),
    85 => (x"99",x"ff",x"c3",x"29"),
    86 => (x"66",x"d0",x"7c",x"71"),
    87 => (x"c3",x"29",x"c8",x"49"),
    88 => (x"7c",x"71",x"99",x"ff"),
    89 => (x"c3",x"49",x"66",x"d0"),
    90 => (x"7c",x"71",x"99",x"ff"),
    91 => (x"29",x"d0",x"49",x"72"),
    92 => (x"71",x"99",x"ff",x"c3"),
    93 => (x"c9",x"4b",x"6c",x"7c"),
    94 => (x"c3",x"4d",x"ff",x"f0"),
    95 => (x"d0",x"05",x"ab",x"ff"),
    96 => (x"7c",x"ff",x"c3",x"87"),
    97 => (x"8d",x"c1",x"4b",x"6c"),
    98 => (x"c3",x"87",x"c6",x"02"),
    99 => (x"f0",x"02",x"ab",x"ff"),
   100 => (x"fe",x"48",x"73",x"87"),
   101 => (x"c0",x"1e",x"87",x"c7"),
   102 => (x"48",x"d4",x"ff",x"49"),
   103 => (x"c1",x"78",x"ff",x"c3"),
   104 => (x"b7",x"c8",x"c3",x"81"),
   105 => (x"87",x"f1",x"04",x"a9"),
   106 => (x"73",x"1e",x"4f",x"26"),
   107 => (x"c4",x"87",x"e7",x"1e"),
   108 => (x"c0",x"4b",x"df",x"f8"),
   109 => (x"f0",x"ff",x"c0",x"1e"),
   110 => (x"fd",x"49",x"f7",x"c1"),
   111 => (x"86",x"c4",x"87",x"e7"),
   112 => (x"c0",x"05",x"a8",x"c1"),
   113 => (x"d4",x"ff",x"87",x"ea"),
   114 => (x"78",x"ff",x"c3",x"48"),
   115 => (x"c0",x"c0",x"c0",x"c1"),
   116 => (x"c0",x"1e",x"c0",x"c0"),
   117 => (x"e9",x"c1",x"f0",x"e1"),
   118 => (x"87",x"c9",x"fd",x"49"),
   119 => (x"98",x"70",x"86",x"c4"),
   120 => (x"ff",x"87",x"ca",x"05"),
   121 => (x"ff",x"c3",x"48",x"d4"),
   122 => (x"cb",x"48",x"c1",x"78"),
   123 => (x"87",x"e6",x"fe",x"87"),
   124 => (x"fe",x"05",x"8b",x"c1"),
   125 => (x"48",x"c0",x"87",x"fd"),
   126 => (x"1e",x"87",x"e6",x"fc"),
   127 => (x"d4",x"ff",x"1e",x"73"),
   128 => (x"78",x"ff",x"c3",x"48"),
   129 => (x"1e",x"c0",x"4b",x"d3"),
   130 => (x"c1",x"f0",x"ff",x"c0"),
   131 => (x"d4",x"fc",x"49",x"c1"),
   132 => (x"70",x"86",x"c4",x"87"),
   133 => (x"87",x"ca",x"05",x"98"),
   134 => (x"c3",x"48",x"d4",x"ff"),
   135 => (x"48",x"c1",x"78",x"ff"),
   136 => (x"f1",x"fd",x"87",x"cb"),
   137 => (x"05",x"8b",x"c1",x"87"),
   138 => (x"c0",x"87",x"db",x"ff"),
   139 => (x"87",x"f1",x"fb",x"48"),
   140 => (x"5c",x"5b",x"5e",x"0e"),
   141 => (x"4c",x"d4",x"ff",x"0e"),
   142 => (x"c6",x"87",x"db",x"fd"),
   143 => (x"e1",x"c0",x"1e",x"ea"),
   144 => (x"49",x"c8",x"c1",x"f0"),
   145 => (x"c4",x"87",x"de",x"fb"),
   146 => (x"02",x"a8",x"c1",x"86"),
   147 => (x"ea",x"fe",x"87",x"c8"),
   148 => (x"c1",x"48",x"c0",x"87"),
   149 => (x"da",x"fa",x"87",x"e2"),
   150 => (x"cf",x"49",x"70",x"87"),
   151 => (x"c6",x"99",x"ff",x"ff"),
   152 => (x"c8",x"02",x"a9",x"ea"),
   153 => (x"87",x"d3",x"fe",x"87"),
   154 => (x"cb",x"c1",x"48",x"c0"),
   155 => (x"7c",x"ff",x"c3",x"87"),
   156 => (x"fc",x"4b",x"f1",x"c0"),
   157 => (x"98",x"70",x"87",x"f4"),
   158 => (x"87",x"eb",x"c0",x"02"),
   159 => (x"ff",x"c0",x"1e",x"c0"),
   160 => (x"49",x"fa",x"c1",x"f0"),
   161 => (x"c4",x"87",x"de",x"fa"),
   162 => (x"05",x"98",x"70",x"86"),
   163 => (x"ff",x"c3",x"87",x"d9"),
   164 => (x"c3",x"49",x"6c",x"7c"),
   165 => (x"7c",x"7c",x"7c",x"ff"),
   166 => (x"99",x"c0",x"c1",x"7c"),
   167 => (x"c1",x"87",x"c4",x"02"),
   168 => (x"c0",x"87",x"d5",x"48"),
   169 => (x"c2",x"87",x"d1",x"48"),
   170 => (x"87",x"c4",x"05",x"ab"),
   171 => (x"87",x"c8",x"48",x"c0"),
   172 => (x"fe",x"05",x"8b",x"c1"),
   173 => (x"48",x"c0",x"87",x"fd"),
   174 => (x"1e",x"87",x"e4",x"f9"),
   175 => (x"dc",x"c2",x"1e",x"73"),
   176 => (x"78",x"c1",x"48",x"e0"),
   177 => (x"d0",x"ff",x"4b",x"c7"),
   178 => (x"fb",x"78",x"c2",x"48"),
   179 => (x"d0",x"ff",x"87",x"c8"),
   180 => (x"c0",x"78",x"c3",x"48"),
   181 => (x"d0",x"e5",x"c0",x"1e"),
   182 => (x"f9",x"49",x"c0",x"c1"),
   183 => (x"86",x"c4",x"87",x"c7"),
   184 => (x"c1",x"05",x"a8",x"c1"),
   185 => (x"ab",x"c2",x"4b",x"87"),
   186 => (x"c0",x"87",x"c5",x"05"),
   187 => (x"87",x"f9",x"c0",x"48"),
   188 => (x"ff",x"05",x"8b",x"c1"),
   189 => (x"f7",x"fc",x"87",x"d0"),
   190 => (x"e4",x"dc",x"c2",x"87"),
   191 => (x"05",x"98",x"70",x"58"),
   192 => (x"1e",x"c1",x"87",x"cd"),
   193 => (x"c1",x"f0",x"ff",x"c0"),
   194 => (x"d8",x"f8",x"49",x"d0"),
   195 => (x"ff",x"86",x"c4",x"87"),
   196 => (x"ff",x"c3",x"48",x"d4"),
   197 => (x"87",x"e0",x"c4",x"78"),
   198 => (x"58",x"e8",x"dc",x"c2"),
   199 => (x"c2",x"48",x"d0",x"ff"),
   200 => (x"48",x"d4",x"ff",x"78"),
   201 => (x"c1",x"78",x"ff",x"c3"),
   202 => (x"87",x"f5",x"f7",x"48"),
   203 => (x"5c",x"5b",x"5e",x"0e"),
   204 => (x"4a",x"71",x"0e",x"5d"),
   205 => (x"ff",x"4d",x"ff",x"c3"),
   206 => (x"7c",x"75",x"4c",x"d4"),
   207 => (x"c4",x"48",x"d0",x"ff"),
   208 => (x"7c",x"75",x"78",x"c3"),
   209 => (x"ff",x"c0",x"1e",x"72"),
   210 => (x"49",x"d8",x"c1",x"f0"),
   211 => (x"c4",x"87",x"d6",x"f7"),
   212 => (x"02",x"98",x"70",x"86"),
   213 => (x"48",x"c0",x"87",x"c5"),
   214 => (x"75",x"87",x"f0",x"c0"),
   215 => (x"7c",x"fe",x"c3",x"7c"),
   216 => (x"d4",x"1e",x"c0",x"c8"),
   217 => (x"dc",x"f5",x"49",x"66"),
   218 => (x"75",x"86",x"c4",x"87"),
   219 => (x"75",x"7c",x"75",x"7c"),
   220 => (x"e0",x"da",x"d8",x"7c"),
   221 => (x"6c",x"7c",x"75",x"4b"),
   222 => (x"c5",x"05",x"99",x"49"),
   223 => (x"05",x"8b",x"c1",x"87"),
   224 => (x"7c",x"75",x"87",x"f3"),
   225 => (x"c2",x"48",x"d0",x"ff"),
   226 => (x"f6",x"48",x"c1",x"78"),
   227 => (x"ff",x"1e",x"87",x"cf"),
   228 => (x"d0",x"ff",x"4a",x"d4"),
   229 => (x"78",x"d1",x"c4",x"48"),
   230 => (x"c1",x"7a",x"ff",x"c3"),
   231 => (x"87",x"f8",x"05",x"89"),
   232 => (x"73",x"1e",x"4f",x"26"),
   233 => (x"c5",x"4b",x"71",x"1e"),
   234 => (x"4a",x"df",x"cd",x"ee"),
   235 => (x"c3",x"48",x"d4",x"ff"),
   236 => (x"48",x"68",x"78",x"ff"),
   237 => (x"02",x"a8",x"fe",x"c3"),
   238 => (x"8a",x"c1",x"87",x"c5"),
   239 => (x"72",x"87",x"ed",x"05"),
   240 => (x"87",x"c5",x"05",x"9a"),
   241 => (x"ea",x"c0",x"48",x"c0"),
   242 => (x"02",x"9b",x"73",x"87"),
   243 => (x"66",x"c8",x"87",x"cc"),
   244 => (x"f4",x"49",x"73",x"1e"),
   245 => (x"86",x"c4",x"87",x"c5"),
   246 => (x"66",x"c8",x"87",x"c6"),
   247 => (x"87",x"ee",x"fe",x"49"),
   248 => (x"c3",x"48",x"d4",x"ff"),
   249 => (x"73",x"78",x"78",x"ff"),
   250 => (x"87",x"c5",x"05",x"9b"),
   251 => (x"d0",x"48",x"d0",x"ff"),
   252 => (x"f4",x"48",x"c1",x"78"),
   253 => (x"73",x"1e",x"87",x"eb"),
   254 => (x"c0",x"4a",x"71",x"1e"),
   255 => (x"48",x"d4",x"ff",x"4b"),
   256 => (x"ff",x"78",x"ff",x"c3"),
   257 => (x"c3",x"c4",x"48",x"d0"),
   258 => (x"48",x"d4",x"ff",x"78"),
   259 => (x"72",x"78",x"ff",x"c3"),
   260 => (x"f0",x"ff",x"c0",x"1e"),
   261 => (x"f4",x"49",x"d1",x"c1"),
   262 => (x"86",x"c4",x"87",x"cb"),
   263 => (x"cd",x"05",x"98",x"70"),
   264 => (x"1e",x"c0",x"c8",x"87"),
   265 => (x"fd",x"49",x"66",x"cc"),
   266 => (x"86",x"c4",x"87",x"f8"),
   267 => (x"d0",x"ff",x"4b",x"70"),
   268 => (x"73",x"78",x"c2",x"48"),
   269 => (x"87",x"e9",x"f3",x"48"),
   270 => (x"5c",x"5b",x"5e",x"0e"),
   271 => (x"1e",x"c0",x"0e",x"5d"),
   272 => (x"c1",x"f0",x"ff",x"c0"),
   273 => (x"dc",x"f3",x"49",x"c9"),
   274 => (x"c2",x"1e",x"d2",x"87"),
   275 => (x"fd",x"49",x"e8",x"dc"),
   276 => (x"86",x"c8",x"87",x"d0"),
   277 => (x"84",x"c1",x"4c",x"c0"),
   278 => (x"04",x"ac",x"b7",x"d2"),
   279 => (x"dc",x"c2",x"87",x"f8"),
   280 => (x"49",x"bf",x"97",x"e8"),
   281 => (x"c1",x"99",x"c0",x"c3"),
   282 => (x"c0",x"05",x"a9",x"c0"),
   283 => (x"dc",x"c2",x"87",x"e7"),
   284 => (x"49",x"bf",x"97",x"ef"),
   285 => (x"dc",x"c2",x"31",x"d0"),
   286 => (x"4a",x"bf",x"97",x"f0"),
   287 => (x"b1",x"72",x"32",x"c8"),
   288 => (x"97",x"f1",x"dc",x"c2"),
   289 => (x"71",x"b1",x"4a",x"bf"),
   290 => (x"ff",x"ff",x"cf",x"4c"),
   291 => (x"84",x"c1",x"9c",x"ff"),
   292 => (x"e7",x"c1",x"34",x"ca"),
   293 => (x"f1",x"dc",x"c2",x"87"),
   294 => (x"c1",x"49",x"bf",x"97"),
   295 => (x"c2",x"99",x"c6",x"31"),
   296 => (x"bf",x"97",x"f2",x"dc"),
   297 => (x"2a",x"b7",x"c7",x"4a"),
   298 => (x"dc",x"c2",x"b1",x"72"),
   299 => (x"4a",x"bf",x"97",x"ed"),
   300 => (x"c2",x"9d",x"cf",x"4d"),
   301 => (x"bf",x"97",x"ee",x"dc"),
   302 => (x"ca",x"9a",x"c3",x"4a"),
   303 => (x"ef",x"dc",x"c2",x"32"),
   304 => (x"c2",x"4b",x"bf",x"97"),
   305 => (x"c2",x"b2",x"73",x"33"),
   306 => (x"bf",x"97",x"f0",x"dc"),
   307 => (x"9b",x"c0",x"c3",x"4b"),
   308 => (x"73",x"2b",x"b7",x"c6"),
   309 => (x"c1",x"81",x"c2",x"b2"),
   310 => (x"70",x"30",x"71",x"48"),
   311 => (x"75",x"48",x"c1",x"49"),
   312 => (x"72",x"4d",x"70",x"30"),
   313 => (x"71",x"84",x"c1",x"4c"),
   314 => (x"b7",x"c0",x"c8",x"94"),
   315 => (x"87",x"cc",x"06",x"ad"),
   316 => (x"2d",x"b7",x"34",x"c1"),
   317 => (x"ad",x"b7",x"c0",x"c8"),
   318 => (x"87",x"f4",x"ff",x"01"),
   319 => (x"dc",x"f0",x"48",x"74"),
   320 => (x"5b",x"5e",x"0e",x"87"),
   321 => (x"f8",x"0e",x"5d",x"5c"),
   322 => (x"ce",x"e5",x"c2",x"86"),
   323 => (x"c2",x"78",x"c0",x"48"),
   324 => (x"c0",x"1e",x"c6",x"dd"),
   325 => (x"87",x"de",x"fb",x"49"),
   326 => (x"98",x"70",x"86",x"c4"),
   327 => (x"c0",x"87",x"c5",x"05"),
   328 => (x"87",x"ce",x"c9",x"48"),
   329 => (x"7e",x"c1",x"4d",x"c0"),
   330 => (x"bf",x"cb",x"f2",x"c0"),
   331 => (x"fc",x"dd",x"c2",x"49"),
   332 => (x"4b",x"c8",x"71",x"4a"),
   333 => (x"70",x"87",x"f3",x"ec"),
   334 => (x"87",x"c2",x"05",x"98"),
   335 => (x"f2",x"c0",x"7e",x"c0"),
   336 => (x"c2",x"49",x"bf",x"c7"),
   337 => (x"71",x"4a",x"d8",x"de"),
   338 => (x"dd",x"ec",x"4b",x"c8"),
   339 => (x"05",x"98",x"70",x"87"),
   340 => (x"7e",x"c0",x"87",x"c2"),
   341 => (x"fd",x"c0",x"02",x"6e"),
   342 => (x"cc",x"e4",x"c2",x"87"),
   343 => (x"e5",x"c2",x"4d",x"bf"),
   344 => (x"7e",x"bf",x"9f",x"c4"),
   345 => (x"ea",x"d6",x"c5",x"48"),
   346 => (x"87",x"c7",x"05",x"a8"),
   347 => (x"bf",x"cc",x"e4",x"c2"),
   348 => (x"6e",x"87",x"ce",x"4d"),
   349 => (x"d5",x"e9",x"ca",x"48"),
   350 => (x"87",x"c5",x"02",x"a8"),
   351 => (x"f1",x"c7",x"48",x"c0"),
   352 => (x"c6",x"dd",x"c2",x"87"),
   353 => (x"f9",x"49",x"75",x"1e"),
   354 => (x"86",x"c4",x"87",x"ec"),
   355 => (x"c5",x"05",x"98",x"70"),
   356 => (x"c7",x"48",x"c0",x"87"),
   357 => (x"f2",x"c0",x"87",x"dc"),
   358 => (x"c2",x"49",x"bf",x"c7"),
   359 => (x"71",x"4a",x"d8",x"de"),
   360 => (x"c5",x"eb",x"4b",x"c8"),
   361 => (x"05",x"98",x"70",x"87"),
   362 => (x"e5",x"c2",x"87",x"c8"),
   363 => (x"78",x"c1",x"48",x"ce"),
   364 => (x"f2",x"c0",x"87",x"da"),
   365 => (x"c2",x"49",x"bf",x"cb"),
   366 => (x"71",x"4a",x"fc",x"dd"),
   367 => (x"e9",x"ea",x"4b",x"c8"),
   368 => (x"02",x"98",x"70",x"87"),
   369 => (x"c0",x"87",x"c5",x"c0"),
   370 => (x"87",x"e6",x"c6",x"48"),
   371 => (x"97",x"c4",x"e5",x"c2"),
   372 => (x"d5",x"c1",x"49",x"bf"),
   373 => (x"cd",x"c0",x"05",x"a9"),
   374 => (x"c5",x"e5",x"c2",x"87"),
   375 => (x"c2",x"49",x"bf",x"97"),
   376 => (x"c0",x"02",x"a9",x"ea"),
   377 => (x"48",x"c0",x"87",x"c5"),
   378 => (x"c2",x"87",x"c7",x"c6"),
   379 => (x"bf",x"97",x"c6",x"dd"),
   380 => (x"e9",x"c3",x"48",x"7e"),
   381 => (x"ce",x"c0",x"02",x"a8"),
   382 => (x"c3",x"48",x"6e",x"87"),
   383 => (x"c0",x"02",x"a8",x"eb"),
   384 => (x"48",x"c0",x"87",x"c5"),
   385 => (x"c2",x"87",x"eb",x"c5"),
   386 => (x"bf",x"97",x"d1",x"dd"),
   387 => (x"c0",x"05",x"99",x"49"),
   388 => (x"dd",x"c2",x"87",x"cc"),
   389 => (x"49",x"bf",x"97",x"d2"),
   390 => (x"c0",x"02",x"a9",x"c2"),
   391 => (x"48",x"c0",x"87",x"c5"),
   392 => (x"c2",x"87",x"cf",x"c5"),
   393 => (x"bf",x"97",x"d3",x"dd"),
   394 => (x"ca",x"e5",x"c2",x"48"),
   395 => (x"48",x"4c",x"70",x"58"),
   396 => (x"e5",x"c2",x"88",x"c1"),
   397 => (x"dd",x"c2",x"58",x"ce"),
   398 => (x"49",x"bf",x"97",x"d4"),
   399 => (x"dd",x"c2",x"81",x"75"),
   400 => (x"4a",x"bf",x"97",x"d5"),
   401 => (x"a1",x"72",x"32",x"c8"),
   402 => (x"db",x"e9",x"c2",x"7e"),
   403 => (x"c2",x"78",x"6e",x"48"),
   404 => (x"bf",x"97",x"d6",x"dd"),
   405 => (x"58",x"a6",x"c8",x"48"),
   406 => (x"bf",x"ce",x"e5",x"c2"),
   407 => (x"87",x"d4",x"c2",x"02"),
   408 => (x"bf",x"c7",x"f2",x"c0"),
   409 => (x"d8",x"de",x"c2",x"49"),
   410 => (x"4b",x"c8",x"71",x"4a"),
   411 => (x"70",x"87",x"fb",x"e7"),
   412 => (x"c5",x"c0",x"02",x"98"),
   413 => (x"c3",x"48",x"c0",x"87"),
   414 => (x"e5",x"c2",x"87",x"f8"),
   415 => (x"c2",x"4c",x"bf",x"c6"),
   416 => (x"c2",x"5c",x"ef",x"e9"),
   417 => (x"bf",x"97",x"eb",x"dd"),
   418 => (x"c2",x"31",x"c8",x"49"),
   419 => (x"bf",x"97",x"ea",x"dd"),
   420 => (x"c2",x"49",x"a1",x"4a"),
   421 => (x"bf",x"97",x"ec",x"dd"),
   422 => (x"72",x"32",x"d0",x"4a"),
   423 => (x"dd",x"c2",x"49",x"a1"),
   424 => (x"4a",x"bf",x"97",x"ed"),
   425 => (x"a1",x"72",x"32",x"d8"),
   426 => (x"91",x"66",x"c4",x"49"),
   427 => (x"bf",x"db",x"e9",x"c2"),
   428 => (x"e3",x"e9",x"c2",x"81"),
   429 => (x"f3",x"dd",x"c2",x"59"),
   430 => (x"c8",x"4a",x"bf",x"97"),
   431 => (x"f2",x"dd",x"c2",x"32"),
   432 => (x"a2",x"4b",x"bf",x"97"),
   433 => (x"f4",x"dd",x"c2",x"4a"),
   434 => (x"d0",x"4b",x"bf",x"97"),
   435 => (x"4a",x"a2",x"73",x"33"),
   436 => (x"97",x"f5",x"dd",x"c2"),
   437 => (x"9b",x"cf",x"4b",x"bf"),
   438 => (x"a2",x"73",x"33",x"d8"),
   439 => (x"e7",x"e9",x"c2",x"4a"),
   440 => (x"e3",x"e9",x"c2",x"5a"),
   441 => (x"8a",x"c2",x"4a",x"bf"),
   442 => (x"e9",x"c2",x"92",x"74"),
   443 => (x"a1",x"72",x"48",x"e7"),
   444 => (x"87",x"ca",x"c1",x"78"),
   445 => (x"97",x"d8",x"dd",x"c2"),
   446 => (x"31",x"c8",x"49",x"bf"),
   447 => (x"97",x"d7",x"dd",x"c2"),
   448 => (x"49",x"a1",x"4a",x"bf"),
   449 => (x"59",x"d6",x"e5",x"c2"),
   450 => (x"bf",x"d2",x"e5",x"c2"),
   451 => (x"c7",x"31",x"c5",x"49"),
   452 => (x"29",x"c9",x"81",x"ff"),
   453 => (x"59",x"ef",x"e9",x"c2"),
   454 => (x"97",x"dd",x"dd",x"c2"),
   455 => (x"32",x"c8",x"4a",x"bf"),
   456 => (x"97",x"dc",x"dd",x"c2"),
   457 => (x"4a",x"a2",x"4b",x"bf"),
   458 => (x"6e",x"92",x"66",x"c4"),
   459 => (x"eb",x"e9",x"c2",x"82"),
   460 => (x"e3",x"e9",x"c2",x"5a"),
   461 => (x"c2",x"78",x"c0",x"48"),
   462 => (x"72",x"48",x"df",x"e9"),
   463 => (x"e9",x"c2",x"78",x"a1"),
   464 => (x"e9",x"c2",x"48",x"ef"),
   465 => (x"c2",x"78",x"bf",x"e3"),
   466 => (x"c2",x"48",x"f3",x"e9"),
   467 => (x"78",x"bf",x"e7",x"e9"),
   468 => (x"bf",x"ce",x"e5",x"c2"),
   469 => (x"87",x"c9",x"c0",x"02"),
   470 => (x"30",x"c4",x"48",x"74"),
   471 => (x"c9",x"c0",x"7e",x"70"),
   472 => (x"eb",x"e9",x"c2",x"87"),
   473 => (x"30",x"c4",x"48",x"bf"),
   474 => (x"e5",x"c2",x"7e",x"70"),
   475 => (x"78",x"6e",x"48",x"d2"),
   476 => (x"8e",x"f8",x"48",x"c1"),
   477 => (x"4c",x"26",x"4d",x"26"),
   478 => (x"4f",x"26",x"4b",x"26"),
   479 => (x"5c",x"5b",x"5e",x"0e"),
   480 => (x"4a",x"71",x"0e",x"5d"),
   481 => (x"bf",x"ce",x"e5",x"c2"),
   482 => (x"72",x"87",x"cb",x"02"),
   483 => (x"72",x"2b",x"c7",x"4b"),
   484 => (x"9c",x"ff",x"c1",x"4c"),
   485 => (x"4b",x"72",x"87",x"c9"),
   486 => (x"4c",x"72",x"2b",x"c8"),
   487 => (x"c2",x"9c",x"ff",x"c3"),
   488 => (x"83",x"bf",x"db",x"e9"),
   489 => (x"bf",x"c3",x"f2",x"c0"),
   490 => (x"87",x"d9",x"02",x"ab"),
   491 => (x"5b",x"c7",x"f2",x"c0"),
   492 => (x"1e",x"c6",x"dd",x"c2"),
   493 => (x"fd",x"f0",x"49",x"73"),
   494 => (x"70",x"86",x"c4",x"87"),
   495 => (x"87",x"c5",x"05",x"98"),
   496 => (x"e6",x"c0",x"48",x"c0"),
   497 => (x"ce",x"e5",x"c2",x"87"),
   498 => (x"87",x"d2",x"02",x"bf"),
   499 => (x"91",x"c4",x"49",x"74"),
   500 => (x"81",x"c6",x"dd",x"c2"),
   501 => (x"ff",x"cf",x"4d",x"69"),
   502 => (x"9d",x"ff",x"ff",x"ff"),
   503 => (x"49",x"74",x"87",x"cb"),
   504 => (x"dd",x"c2",x"91",x"c2"),
   505 => (x"69",x"9f",x"81",x"c6"),
   506 => (x"fe",x"48",x"75",x"4d"),
   507 => (x"5e",x"0e",x"87",x"c6"),
   508 => (x"0e",x"5d",x"5c",x"5b"),
   509 => (x"c0",x"4d",x"71",x"1e"),
   510 => (x"ca",x"49",x"c1",x"1e"),
   511 => (x"86",x"c4",x"87",x"ee"),
   512 => (x"02",x"9c",x"4c",x"70"),
   513 => (x"c2",x"87",x"c0",x"c1"),
   514 => (x"75",x"4a",x"d6",x"e5"),
   515 => (x"87",x"ff",x"e0",x"49"),
   516 => (x"c0",x"02",x"98",x"70"),
   517 => (x"4a",x"74",x"87",x"f1"),
   518 => (x"4b",x"cb",x"49",x"75"),
   519 => (x"70",x"87",x"e5",x"e1"),
   520 => (x"e2",x"c0",x"02",x"98"),
   521 => (x"74",x"1e",x"c0",x"87"),
   522 => (x"87",x"c7",x"02",x"9c"),
   523 => (x"c0",x"48",x"a6",x"c4"),
   524 => (x"c4",x"87",x"c5",x"78"),
   525 => (x"78",x"c1",x"48",x"a6"),
   526 => (x"c9",x"49",x"66",x"c4"),
   527 => (x"86",x"c4",x"87",x"ee"),
   528 => (x"05",x"9c",x"4c",x"70"),
   529 => (x"74",x"87",x"c0",x"ff"),
   530 => (x"e7",x"fc",x"26",x"48"),
   531 => (x"5b",x"5e",x"0e",x"87"),
   532 => (x"1e",x"0e",x"5d",x"5c"),
   533 => (x"05",x"9b",x"4b",x"71"),
   534 => (x"48",x"c0",x"87",x"c5"),
   535 => (x"c8",x"87",x"e5",x"c1"),
   536 => (x"7d",x"c0",x"4d",x"a3"),
   537 => (x"c7",x"02",x"66",x"d4"),
   538 => (x"97",x"66",x"d4",x"87"),
   539 => (x"87",x"c5",x"05",x"bf"),
   540 => (x"cf",x"c1",x"48",x"c0"),
   541 => (x"49",x"66",x"d4",x"87"),
   542 => (x"70",x"87",x"f3",x"fd"),
   543 => (x"c1",x"02",x"9c",x"4c"),
   544 => (x"a4",x"dc",x"87",x"c0"),
   545 => (x"da",x"7d",x"69",x"49"),
   546 => (x"a3",x"c4",x"49",x"a4"),
   547 => (x"7a",x"69",x"9f",x"4a"),
   548 => (x"bf",x"ce",x"e5",x"c2"),
   549 => (x"d4",x"87",x"d2",x"02"),
   550 => (x"69",x"9f",x"49",x"a4"),
   551 => (x"ff",x"ff",x"c0",x"49"),
   552 => (x"d0",x"48",x"71",x"99"),
   553 => (x"c2",x"7e",x"70",x"30"),
   554 => (x"6e",x"7e",x"c0",x"87"),
   555 => (x"80",x"6a",x"48",x"49"),
   556 => (x"7b",x"c0",x"7a",x"70"),
   557 => (x"6a",x"49",x"a3",x"cc"),
   558 => (x"49",x"a3",x"d0",x"79"),
   559 => (x"48",x"74",x"79",x"c0"),
   560 => (x"48",x"c0",x"87",x"c2"),
   561 => (x"87",x"ec",x"fa",x"26"),
   562 => (x"5c",x"5b",x"5e",x"0e"),
   563 => (x"4c",x"71",x"0e",x"5d"),
   564 => (x"48",x"c3",x"f2",x"c0"),
   565 => (x"9c",x"74",x"78",x"ff"),
   566 => (x"87",x"ca",x"c1",x"02"),
   567 => (x"69",x"49",x"a4",x"c8"),
   568 => (x"87",x"c2",x"c1",x"02"),
   569 => (x"6c",x"4a",x"66",x"d0"),
   570 => (x"a6",x"d4",x"82",x"49"),
   571 => (x"4d",x"66",x"d0",x"5a"),
   572 => (x"ca",x"e5",x"c2",x"b9"),
   573 => (x"ba",x"ff",x"4a",x"bf"),
   574 => (x"99",x"71",x"99",x"72"),
   575 => (x"87",x"e4",x"c0",x"02"),
   576 => (x"6b",x"4b",x"a4",x"c4"),
   577 => (x"87",x"f4",x"f9",x"49"),
   578 => (x"e5",x"c2",x"7b",x"70"),
   579 => (x"6c",x"49",x"bf",x"c6"),
   580 => (x"75",x"7c",x"71",x"81"),
   581 => (x"ca",x"e5",x"c2",x"b9"),
   582 => (x"ba",x"ff",x"4a",x"bf"),
   583 => (x"99",x"71",x"99",x"72"),
   584 => (x"87",x"dc",x"ff",x"05"),
   585 => (x"cb",x"f9",x"7c",x"75"),
   586 => (x"1e",x"73",x"1e",x"87"),
   587 => (x"02",x"9b",x"4b",x"71"),
   588 => (x"a3",x"c8",x"87",x"c7"),
   589 => (x"c5",x"05",x"69",x"49"),
   590 => (x"c0",x"48",x"c0",x"87"),
   591 => (x"e9",x"c2",x"87",x"eb"),
   592 => (x"c4",x"4a",x"bf",x"df"),
   593 => (x"49",x"69",x"49",x"a3"),
   594 => (x"e5",x"c2",x"89",x"c2"),
   595 => (x"71",x"91",x"bf",x"c6"),
   596 => (x"e5",x"c2",x"4a",x"a2"),
   597 => (x"6b",x"49",x"bf",x"ca"),
   598 => (x"4a",x"a2",x"71",x"99"),
   599 => (x"72",x"1e",x"66",x"c8"),
   600 => (x"87",x"d2",x"ea",x"49"),
   601 => (x"49",x"70",x"86",x"c4"),
   602 => (x"87",x"cc",x"f8",x"48"),
   603 => (x"71",x"1e",x"73",x"1e"),
   604 => (x"c7",x"02",x"9b",x"4b"),
   605 => (x"49",x"a3",x"c8",x"87"),
   606 => (x"87",x"c5",x"05",x"69"),
   607 => (x"eb",x"c0",x"48",x"c0"),
   608 => (x"df",x"e9",x"c2",x"87"),
   609 => (x"a3",x"c4",x"4a",x"bf"),
   610 => (x"c2",x"49",x"69",x"49"),
   611 => (x"c6",x"e5",x"c2",x"89"),
   612 => (x"a2",x"71",x"91",x"bf"),
   613 => (x"ca",x"e5",x"c2",x"4a"),
   614 => (x"99",x"6b",x"49",x"bf"),
   615 => (x"c8",x"4a",x"a2",x"71"),
   616 => (x"49",x"72",x"1e",x"66"),
   617 => (x"c4",x"87",x"c5",x"e6"),
   618 => (x"48",x"49",x"70",x"86"),
   619 => (x"0e",x"87",x"c9",x"f7"),
   620 => (x"5d",x"5c",x"5b",x"5e"),
   621 => (x"4b",x"71",x"1e",x"0e"),
   622 => (x"c9",x"4c",x"66",x"d4"),
   623 => (x"02",x"9b",x"73",x"2c"),
   624 => (x"c8",x"87",x"cf",x"c1"),
   625 => (x"02",x"69",x"49",x"a3"),
   626 => (x"d0",x"87",x"c7",x"c1"),
   627 => (x"66",x"d4",x"4d",x"a3"),
   628 => (x"ca",x"e5",x"c2",x"7d"),
   629 => (x"b9",x"ff",x"49",x"bf"),
   630 => (x"7e",x"99",x"4a",x"6b"),
   631 => (x"cd",x"03",x"ac",x"71"),
   632 => (x"7d",x"7b",x"c0",x"87"),
   633 => (x"c4",x"4a",x"a3",x"cc"),
   634 => (x"79",x"6a",x"49",x"a3"),
   635 => (x"8c",x"72",x"87",x"c2"),
   636 => (x"dd",x"02",x"9c",x"74"),
   637 => (x"73",x"1e",x"49",x"87"),
   638 => (x"87",x"cc",x"fb",x"49"),
   639 => (x"66",x"d4",x"86",x"c4"),
   640 => (x"99",x"ff",x"c7",x"49"),
   641 => (x"c2",x"87",x"cb",x"02"),
   642 => (x"73",x"1e",x"c6",x"dd"),
   643 => (x"87",x"d9",x"fc",x"49"),
   644 => (x"f5",x"26",x"86",x"c4"),
   645 => (x"73",x"1e",x"87",x"de"),
   646 => (x"9b",x"4b",x"71",x"1e"),
   647 => (x"87",x"e4",x"c0",x"02"),
   648 => (x"5b",x"f3",x"e9",x"c2"),
   649 => (x"8a",x"c2",x"4a",x"73"),
   650 => (x"bf",x"c6",x"e5",x"c2"),
   651 => (x"e9",x"c2",x"92",x"49"),
   652 => (x"72",x"48",x"bf",x"df"),
   653 => (x"f7",x"e9",x"c2",x"80"),
   654 => (x"c4",x"48",x"71",x"58"),
   655 => (x"d6",x"e5",x"c2",x"30"),
   656 => (x"87",x"ed",x"c0",x"58"),
   657 => (x"48",x"ef",x"e9",x"c2"),
   658 => (x"bf",x"e3",x"e9",x"c2"),
   659 => (x"f3",x"e9",x"c2",x"78"),
   660 => (x"e7",x"e9",x"c2",x"48"),
   661 => (x"e5",x"c2",x"78",x"bf"),
   662 => (x"c9",x"02",x"bf",x"ce"),
   663 => (x"c6",x"e5",x"c2",x"87"),
   664 => (x"31",x"c4",x"49",x"bf"),
   665 => (x"e9",x"c2",x"87",x"c7"),
   666 => (x"c4",x"49",x"bf",x"eb"),
   667 => (x"d6",x"e5",x"c2",x"31"),
   668 => (x"87",x"c4",x"f4",x"59"),
   669 => (x"5c",x"5b",x"5e",x"0e"),
   670 => (x"c0",x"4a",x"71",x"0e"),
   671 => (x"02",x"9a",x"72",x"4b"),
   672 => (x"da",x"87",x"e1",x"c0"),
   673 => (x"69",x"9f",x"49",x"a2"),
   674 => (x"ce",x"e5",x"c2",x"4b"),
   675 => (x"87",x"cf",x"02",x"bf"),
   676 => (x"9f",x"49",x"a2",x"d4"),
   677 => (x"c0",x"4c",x"49",x"69"),
   678 => (x"d0",x"9c",x"ff",x"ff"),
   679 => (x"c0",x"87",x"c2",x"34"),
   680 => (x"b3",x"49",x"74",x"4c"),
   681 => (x"ed",x"fd",x"49",x"73"),
   682 => (x"87",x"ca",x"f3",x"87"),
   683 => (x"5c",x"5b",x"5e",x"0e"),
   684 => (x"86",x"f4",x"0e",x"5d"),
   685 => (x"7e",x"c0",x"4a",x"71"),
   686 => (x"d8",x"02",x"9a",x"72"),
   687 => (x"c2",x"dd",x"c2",x"87"),
   688 => (x"c2",x"78",x"c0",x"48"),
   689 => (x"c2",x"48",x"fa",x"dc"),
   690 => (x"78",x"bf",x"f3",x"e9"),
   691 => (x"48",x"fe",x"dc",x"c2"),
   692 => (x"bf",x"ef",x"e9",x"c2"),
   693 => (x"e3",x"e5",x"c2",x"78"),
   694 => (x"c2",x"50",x"c0",x"48"),
   695 => (x"49",x"bf",x"d2",x"e5"),
   696 => (x"bf",x"c2",x"dd",x"c2"),
   697 => (x"03",x"aa",x"71",x"4a"),
   698 => (x"72",x"87",x"ff",x"c3"),
   699 => (x"05",x"99",x"cf",x"49"),
   700 => (x"c2",x"87",x"e0",x"c0"),
   701 => (x"c2",x"1e",x"c6",x"dd"),
   702 => (x"49",x"bf",x"fa",x"dc"),
   703 => (x"48",x"fa",x"dc",x"c2"),
   704 => (x"71",x"78",x"a1",x"c1"),
   705 => (x"c4",x"87",x"ef",x"e3"),
   706 => (x"ff",x"f1",x"c0",x"86"),
   707 => (x"c6",x"dd",x"c2",x"48"),
   708 => (x"c0",x"87",x"cc",x"78"),
   709 => (x"48",x"bf",x"ff",x"f1"),
   710 => (x"c0",x"80",x"e0",x"c0"),
   711 => (x"c2",x"58",x"c3",x"f2"),
   712 => (x"48",x"bf",x"c2",x"dd"),
   713 => (x"dd",x"c2",x"80",x"c1"),
   714 => (x"7f",x"27",x"58",x"c6"),
   715 => (x"bf",x"00",x"00",x"0c"),
   716 => (x"9d",x"4d",x"bf",x"97"),
   717 => (x"87",x"e2",x"c2",x"02"),
   718 => (x"02",x"ad",x"e5",x"c3"),
   719 => (x"c0",x"87",x"db",x"c2"),
   720 => (x"4b",x"bf",x"ff",x"f1"),
   721 => (x"11",x"49",x"a3",x"cb"),
   722 => (x"05",x"ac",x"cf",x"4c"),
   723 => (x"75",x"87",x"d2",x"c1"),
   724 => (x"c1",x"99",x"df",x"49"),
   725 => (x"c2",x"91",x"cd",x"89"),
   726 => (x"c1",x"81",x"d6",x"e5"),
   727 => (x"51",x"12",x"4a",x"a3"),
   728 => (x"12",x"4a",x"a3",x"c3"),
   729 => (x"4a",x"a3",x"c5",x"51"),
   730 => (x"a3",x"c7",x"51",x"12"),
   731 => (x"c9",x"51",x"12",x"4a"),
   732 => (x"51",x"12",x"4a",x"a3"),
   733 => (x"12",x"4a",x"a3",x"ce"),
   734 => (x"4a",x"a3",x"d0",x"51"),
   735 => (x"a3",x"d2",x"51",x"12"),
   736 => (x"d4",x"51",x"12",x"4a"),
   737 => (x"51",x"12",x"4a",x"a3"),
   738 => (x"12",x"4a",x"a3",x"d6"),
   739 => (x"4a",x"a3",x"d8",x"51"),
   740 => (x"a3",x"dc",x"51",x"12"),
   741 => (x"de",x"51",x"12",x"4a"),
   742 => (x"51",x"12",x"4a",x"a3"),
   743 => (x"f9",x"c0",x"7e",x"c1"),
   744 => (x"c8",x"49",x"74",x"87"),
   745 => (x"ea",x"c0",x"05",x"99"),
   746 => (x"d0",x"49",x"74",x"87"),
   747 => (x"87",x"d0",x"05",x"99"),
   748 => (x"c0",x"02",x"66",x"dc"),
   749 => (x"49",x"73",x"87",x"ca"),
   750 => (x"70",x"0f",x"66",x"dc"),
   751 => (x"87",x"d3",x"02",x"98"),
   752 => (x"c6",x"c0",x"05",x"6e"),
   753 => (x"d6",x"e5",x"c2",x"87"),
   754 => (x"c0",x"50",x"c0",x"48"),
   755 => (x"48",x"bf",x"ff",x"f1"),
   756 => (x"c2",x"87",x"e7",x"c2"),
   757 => (x"c0",x"48",x"e3",x"e5"),
   758 => (x"e5",x"c2",x"7e",x"50"),
   759 => (x"c2",x"49",x"bf",x"d2"),
   760 => (x"4a",x"bf",x"c2",x"dd"),
   761 => (x"fc",x"04",x"aa",x"71"),
   762 => (x"e9",x"c2",x"87",x"c1"),
   763 => (x"c0",x"05",x"bf",x"f3"),
   764 => (x"e5",x"c2",x"87",x"c8"),
   765 => (x"c1",x"02",x"bf",x"ce"),
   766 => (x"f2",x"c0",x"87",x"fe"),
   767 => (x"78",x"ff",x"48",x"c3"),
   768 => (x"bf",x"fe",x"dc",x"c2"),
   769 => (x"87",x"f4",x"ed",x"49"),
   770 => (x"dd",x"c2",x"49",x"70"),
   771 => (x"a6",x"c4",x"59",x"c2"),
   772 => (x"fe",x"dc",x"c2",x"48"),
   773 => (x"e5",x"c2",x"78",x"bf"),
   774 => (x"c0",x"02",x"bf",x"ce"),
   775 => (x"66",x"c4",x"87",x"d8"),
   776 => (x"ff",x"ff",x"cf",x"49"),
   777 => (x"a9",x"99",x"f8",x"ff"),
   778 => (x"87",x"c5",x"c0",x"02"),
   779 => (x"e1",x"c0",x"4d",x"c0"),
   780 => (x"c0",x"4d",x"c1",x"87"),
   781 => (x"66",x"c4",x"87",x"dc"),
   782 => (x"f8",x"ff",x"cf",x"49"),
   783 => (x"c0",x"02",x"a9",x"99"),
   784 => (x"a6",x"c8",x"87",x"c8"),
   785 => (x"c0",x"78",x"c0",x"48"),
   786 => (x"a6",x"c8",x"87",x"c5"),
   787 => (x"c8",x"78",x"c1",x"48"),
   788 => (x"9d",x"75",x"4d",x"66"),
   789 => (x"87",x"e0",x"c0",x"05"),
   790 => (x"c2",x"49",x"66",x"c4"),
   791 => (x"c6",x"e5",x"c2",x"89"),
   792 => (x"c2",x"91",x"4a",x"bf"),
   793 => (x"4a",x"bf",x"df",x"e9"),
   794 => (x"48",x"fa",x"dc",x"c2"),
   795 => (x"c2",x"78",x"a1",x"72"),
   796 => (x"c0",x"48",x"c2",x"dd"),
   797 => (x"87",x"e3",x"f9",x"78"),
   798 => (x"8e",x"f4",x"48",x"c0"),
   799 => (x"00",x"87",x"f5",x"eb"),
   800 => (x"ff",x"00",x"00",x"00"),
   801 => (x"8f",x"ff",x"ff",x"ff"),
   802 => (x"98",x"00",x"00",x"0c"),
   803 => (x"46",x"00",x"00",x"0c"),
   804 => (x"32",x"33",x"54",x"41"),
   805 => (x"00",x"20",x"20",x"20"),
   806 => (x"31",x"54",x"41",x"46"),
   807 => (x"20",x"20",x"20",x"36"),
   808 => (x"d4",x"ff",x"1e",x"00"),
   809 => (x"78",x"ff",x"c3",x"48"),
   810 => (x"4f",x"26",x"48",x"68"),
   811 => (x"48",x"d4",x"ff",x"1e"),
   812 => (x"ff",x"78",x"ff",x"c3"),
   813 => (x"e1",x"c8",x"48",x"d0"),
   814 => (x"48",x"d4",x"ff",x"78"),
   815 => (x"e9",x"c2",x"78",x"d4"),
   816 => (x"d4",x"ff",x"48",x"f7"),
   817 => (x"4f",x"26",x"50",x"bf"),
   818 => (x"48",x"d0",x"ff",x"1e"),
   819 => (x"26",x"78",x"e0",x"c0"),
   820 => (x"cc",x"ff",x"1e",x"4f"),
   821 => (x"99",x"49",x"70",x"87"),
   822 => (x"c0",x"87",x"c6",x"02"),
   823 => (x"f1",x"05",x"a9",x"fb"),
   824 => (x"26",x"48",x"71",x"87"),
   825 => (x"5b",x"5e",x"0e",x"4f"),
   826 => (x"4b",x"71",x"0e",x"5c"),
   827 => (x"f0",x"fe",x"4c",x"c0"),
   828 => (x"99",x"49",x"70",x"87"),
   829 => (x"87",x"f9",x"c0",x"02"),
   830 => (x"02",x"a9",x"ec",x"c0"),
   831 => (x"c0",x"87",x"f2",x"c0"),
   832 => (x"c0",x"02",x"a9",x"fb"),
   833 => (x"66",x"cc",x"87",x"eb"),
   834 => (x"c7",x"03",x"ac",x"b7"),
   835 => (x"02",x"66",x"d0",x"87"),
   836 => (x"53",x"71",x"87",x"c2"),
   837 => (x"c2",x"02",x"99",x"71"),
   838 => (x"fe",x"84",x"c1",x"87"),
   839 => (x"49",x"70",x"87",x"c3"),
   840 => (x"87",x"cd",x"02",x"99"),
   841 => (x"02",x"a9",x"ec",x"c0"),
   842 => (x"fb",x"c0",x"87",x"c7"),
   843 => (x"d5",x"ff",x"05",x"a9"),
   844 => (x"02",x"66",x"d0",x"87"),
   845 => (x"97",x"c0",x"87",x"c3"),
   846 => (x"a9",x"ec",x"c0",x"7b"),
   847 => (x"74",x"87",x"c4",x"05"),
   848 => (x"74",x"87",x"c5",x"4a"),
   849 => (x"8a",x"0a",x"c0",x"4a"),
   850 => (x"87",x"c2",x"48",x"72"),
   851 => (x"4c",x"26",x"4d",x"26"),
   852 => (x"4f",x"26",x"4b",x"26"),
   853 => (x"87",x"c9",x"fd",x"1e"),
   854 => (x"f0",x"c0",x"49",x"70"),
   855 => (x"ca",x"04",x"a9",x"b7"),
   856 => (x"b7",x"f9",x"c0",x"87"),
   857 => (x"87",x"c3",x"01",x"a9"),
   858 => (x"c1",x"89",x"f0",x"c0"),
   859 => (x"04",x"a9",x"b7",x"c1"),
   860 => (x"da",x"c1",x"87",x"ca"),
   861 => (x"c3",x"01",x"a9",x"b7"),
   862 => (x"89",x"f7",x"c0",x"87"),
   863 => (x"4f",x"26",x"48",x"71"),
   864 => (x"5c",x"5b",x"5e",x"0e"),
   865 => (x"ff",x"4a",x"71",x"0e"),
   866 => (x"49",x"72",x"4c",x"d4"),
   867 => (x"70",x"87",x"ea",x"c0"),
   868 => (x"c2",x"02",x"9b",x"4b"),
   869 => (x"ff",x"8b",x"c1",x"87"),
   870 => (x"c5",x"c8",x"48",x"d0"),
   871 => (x"7c",x"d5",x"c1",x"78"),
   872 => (x"31",x"c6",x"49",x"73"),
   873 => (x"97",x"cd",x"db",x"c2"),
   874 => (x"71",x"48",x"4a",x"bf"),
   875 => (x"ff",x"7c",x"70",x"b0"),
   876 => (x"78",x"c4",x"48",x"d0"),
   877 => (x"d5",x"fe",x"48",x"73"),
   878 => (x"5b",x"5e",x"0e",x"87"),
   879 => (x"f8",x"0e",x"5d",x"5c"),
   880 => (x"c0",x"4c",x"71",x"86"),
   881 => (x"87",x"e4",x"fb",x"7e"),
   882 => (x"f9",x"c0",x"4b",x"c0"),
   883 => (x"49",x"bf",x"97",x"e6"),
   884 => (x"cf",x"04",x"a9",x"c0"),
   885 => (x"87",x"f9",x"fb",x"87"),
   886 => (x"f9",x"c0",x"83",x"c1"),
   887 => (x"49",x"bf",x"97",x"e6"),
   888 => (x"87",x"f1",x"06",x"ab"),
   889 => (x"97",x"e6",x"f9",x"c0"),
   890 => (x"87",x"cf",x"02",x"bf"),
   891 => (x"70",x"87",x"f2",x"fa"),
   892 => (x"c6",x"02",x"99",x"49"),
   893 => (x"a9",x"ec",x"c0",x"87"),
   894 => (x"c0",x"87",x"f1",x"05"),
   895 => (x"87",x"e1",x"fa",x"4b"),
   896 => (x"dc",x"fa",x"4d",x"70"),
   897 => (x"58",x"a6",x"c8",x"87"),
   898 => (x"70",x"87",x"d6",x"fa"),
   899 => (x"c8",x"83",x"c1",x"4a"),
   900 => (x"69",x"97",x"49",x"a4"),
   901 => (x"c7",x"02",x"ad",x"49"),
   902 => (x"ad",x"ff",x"c0",x"87"),
   903 => (x"87",x"e7",x"c0",x"05"),
   904 => (x"97",x"49",x"a4",x"c9"),
   905 => (x"66",x"c4",x"49",x"69"),
   906 => (x"87",x"c7",x"02",x"a9"),
   907 => (x"a8",x"ff",x"c0",x"48"),
   908 => (x"ca",x"87",x"d4",x"05"),
   909 => (x"69",x"97",x"49",x"a4"),
   910 => (x"c6",x"02",x"aa",x"49"),
   911 => (x"aa",x"ff",x"c0",x"87"),
   912 => (x"c1",x"87",x"c4",x"05"),
   913 => (x"c0",x"87",x"d0",x"7e"),
   914 => (x"c6",x"02",x"ad",x"ec"),
   915 => (x"ad",x"fb",x"c0",x"87"),
   916 => (x"c0",x"87",x"c4",x"05"),
   917 => (x"6e",x"7e",x"c1",x"4b"),
   918 => (x"87",x"e1",x"fe",x"02"),
   919 => (x"73",x"87",x"e9",x"f9"),
   920 => (x"fb",x"8e",x"f8",x"48"),
   921 => (x"0e",x"00",x"87",x"e6"),
   922 => (x"5d",x"5c",x"5b",x"5e"),
   923 => (x"4b",x"71",x"1e",x"0e"),
   924 => (x"ab",x"4d",x"4c",x"c0"),
   925 => (x"87",x"e8",x"c0",x"04"),
   926 => (x"1e",x"f9",x"f6",x"c0"),
   927 => (x"c4",x"02",x"9d",x"75"),
   928 => (x"c2",x"4a",x"c0",x"87"),
   929 => (x"72",x"4a",x"c1",x"87"),
   930 => (x"87",x"e0",x"f0",x"49"),
   931 => (x"7e",x"70",x"86",x"c4"),
   932 => (x"05",x"6e",x"84",x"c1"),
   933 => (x"4c",x"73",x"87",x"c2"),
   934 => (x"ac",x"73",x"85",x"c1"),
   935 => (x"87",x"d8",x"ff",x"06"),
   936 => (x"26",x"26",x"48",x"6e"),
   937 => (x"26",x"4c",x"26",x"4d"),
   938 => (x"0e",x"4f",x"26",x"4b"),
   939 => (x"5d",x"5c",x"5b",x"5e"),
   940 => (x"4c",x"71",x"1e",x"0e"),
   941 => (x"c2",x"91",x"de",x"49"),
   942 => (x"71",x"4d",x"d1",x"ea"),
   943 => (x"02",x"6d",x"97",x"85"),
   944 => (x"c2",x"87",x"dd",x"c1"),
   945 => (x"4a",x"bf",x"fc",x"e9"),
   946 => (x"49",x"72",x"82",x"74"),
   947 => (x"70",x"87",x"d8",x"fe"),
   948 => (x"c0",x"02",x"6e",x"7e"),
   949 => (x"ea",x"c2",x"87",x"f3"),
   950 => (x"4a",x"6e",x"4b",x"c4"),
   951 => (x"c7",x"ff",x"49",x"cb"),
   952 => (x"4b",x"74",x"87",x"c6"),
   953 => (x"dd",x"c1",x"93",x"cb"),
   954 => (x"83",x"c4",x"83",x"c5"),
   955 => (x"7b",x"e4",x"fc",x"c0"),
   956 => (x"c2",x"c1",x"49",x"74"),
   957 => (x"7b",x"75",x"87",x"fe"),
   958 => (x"97",x"d0",x"ea",x"c2"),
   959 => (x"c2",x"1e",x"49",x"bf"),
   960 => (x"c1",x"49",x"c4",x"ea"),
   961 => (x"c4",x"87",x"c8",x"de"),
   962 => (x"c1",x"49",x"74",x"86"),
   963 => (x"c0",x"87",x"e5",x"c2"),
   964 => (x"c4",x"c4",x"c1",x"49"),
   965 => (x"f8",x"e9",x"c2",x"87"),
   966 => (x"c1",x"78",x"c0",x"48"),
   967 => (x"87",x"f9",x"dc",x"49"),
   968 => (x"87",x"ff",x"fd",x"26"),
   969 => (x"64",x"61",x"6f",x"4c"),
   970 => (x"2e",x"67",x"6e",x"69"),
   971 => (x"0e",x"00",x"2e",x"2e"),
   972 => (x"0e",x"5c",x"5b",x"5e"),
   973 => (x"c2",x"4a",x"4b",x"71"),
   974 => (x"82",x"bf",x"fc",x"e9"),
   975 => (x"e6",x"fc",x"49",x"72"),
   976 => (x"9c",x"4c",x"70",x"87"),
   977 => (x"49",x"87",x"c4",x"02"),
   978 => (x"c2",x"87",x"e9",x"ec"),
   979 => (x"c0",x"48",x"fc",x"e9"),
   980 => (x"dc",x"49",x"c1",x"78"),
   981 => (x"cc",x"fd",x"87",x"c3"),
   982 => (x"5b",x"5e",x"0e",x"87"),
   983 => (x"f4",x"0e",x"5d",x"5c"),
   984 => (x"c6",x"dd",x"c2",x"86"),
   985 => (x"c4",x"4c",x"c0",x"4d"),
   986 => (x"78",x"c0",x"48",x"a6"),
   987 => (x"bf",x"fc",x"e9",x"c2"),
   988 => (x"06",x"a9",x"c0",x"49"),
   989 => (x"c2",x"87",x"c1",x"c1"),
   990 => (x"98",x"48",x"c6",x"dd"),
   991 => (x"87",x"f8",x"c0",x"02"),
   992 => (x"1e",x"f9",x"f6",x"c0"),
   993 => (x"c7",x"02",x"66",x"c8"),
   994 => (x"48",x"a6",x"c4",x"87"),
   995 => (x"87",x"c5",x"78",x"c0"),
   996 => (x"c1",x"48",x"a6",x"c4"),
   997 => (x"49",x"66",x"c4",x"78"),
   998 => (x"c4",x"87",x"d1",x"ec"),
   999 => (x"c1",x"4d",x"70",x"86"),
  1000 => (x"48",x"66",x"c4",x"84"),
  1001 => (x"a6",x"c8",x"80",x"c1"),
  1002 => (x"fc",x"e9",x"c2",x"58"),
  1003 => (x"03",x"ac",x"49",x"bf"),
  1004 => (x"9d",x"75",x"87",x"c6"),
  1005 => (x"87",x"c8",x"ff",x"05"),
  1006 => (x"9d",x"75",x"4c",x"c0"),
  1007 => (x"87",x"e0",x"c3",x"02"),
  1008 => (x"1e",x"f9",x"f6",x"c0"),
  1009 => (x"c7",x"02",x"66",x"c8"),
  1010 => (x"48",x"a6",x"cc",x"87"),
  1011 => (x"87",x"c5",x"78",x"c0"),
  1012 => (x"c1",x"48",x"a6",x"cc"),
  1013 => (x"49",x"66",x"cc",x"78"),
  1014 => (x"c4",x"87",x"d1",x"eb"),
  1015 => (x"6e",x"7e",x"70",x"86"),
  1016 => (x"87",x"e9",x"c2",x"02"),
  1017 => (x"81",x"cb",x"49",x"6e"),
  1018 => (x"d0",x"49",x"69",x"97"),
  1019 => (x"d6",x"c1",x"02",x"99"),
  1020 => (x"ef",x"fc",x"c0",x"87"),
  1021 => (x"cb",x"49",x"74",x"4a"),
  1022 => (x"c5",x"dd",x"c1",x"91"),
  1023 => (x"c8",x"79",x"72",x"81"),
  1024 => (x"51",x"ff",x"c3",x"81"),
  1025 => (x"91",x"de",x"49",x"74"),
  1026 => (x"4d",x"d1",x"ea",x"c2"),
  1027 => (x"c1",x"c2",x"85",x"71"),
  1028 => (x"a5",x"c1",x"7d",x"97"),
  1029 => (x"51",x"e0",x"c0",x"49"),
  1030 => (x"97",x"d6",x"e5",x"c2"),
  1031 => (x"87",x"d2",x"02",x"bf"),
  1032 => (x"a5",x"c2",x"84",x"c1"),
  1033 => (x"d6",x"e5",x"c2",x"4b"),
  1034 => (x"ff",x"49",x"db",x"4a"),
  1035 => (x"c1",x"87",x"f9",x"c1"),
  1036 => (x"a5",x"cd",x"87",x"db"),
  1037 => (x"c1",x"51",x"c0",x"49"),
  1038 => (x"4b",x"a5",x"c2",x"84"),
  1039 => (x"49",x"cb",x"4a",x"6e"),
  1040 => (x"87",x"e4",x"c1",x"ff"),
  1041 => (x"c0",x"87",x"c6",x"c1"),
  1042 => (x"74",x"4a",x"eb",x"fa"),
  1043 => (x"c1",x"91",x"cb",x"49"),
  1044 => (x"72",x"81",x"c5",x"dd"),
  1045 => (x"d6",x"e5",x"c2",x"79"),
  1046 => (x"d8",x"02",x"bf",x"97"),
  1047 => (x"de",x"49",x"74",x"87"),
  1048 => (x"c2",x"84",x"c1",x"91"),
  1049 => (x"71",x"4b",x"d1",x"ea"),
  1050 => (x"d6",x"e5",x"c2",x"83"),
  1051 => (x"ff",x"49",x"dd",x"4a"),
  1052 => (x"d8",x"87",x"f5",x"c0"),
  1053 => (x"de",x"4b",x"74",x"87"),
  1054 => (x"d1",x"ea",x"c2",x"93"),
  1055 => (x"49",x"a3",x"cb",x"83"),
  1056 => (x"84",x"c1",x"51",x"c0"),
  1057 => (x"cb",x"4a",x"6e",x"73"),
  1058 => (x"db",x"c0",x"ff",x"49"),
  1059 => (x"48",x"66",x"c4",x"87"),
  1060 => (x"a6",x"c8",x"80",x"c1"),
  1061 => (x"03",x"ac",x"c7",x"58"),
  1062 => (x"6e",x"87",x"c5",x"c0"),
  1063 => (x"87",x"e0",x"fc",x"05"),
  1064 => (x"8e",x"f4",x"48",x"74"),
  1065 => (x"1e",x"87",x"fc",x"f7"),
  1066 => (x"4b",x"71",x"1e",x"73"),
  1067 => (x"c1",x"91",x"cb",x"49"),
  1068 => (x"c8",x"81",x"c5",x"dd"),
  1069 => (x"db",x"c2",x"4a",x"a1"),
  1070 => (x"50",x"12",x"48",x"cd"),
  1071 => (x"c0",x"4a",x"a1",x"c9"),
  1072 => (x"12",x"48",x"e6",x"f9"),
  1073 => (x"c2",x"81",x"ca",x"50"),
  1074 => (x"11",x"48",x"d0",x"ea"),
  1075 => (x"d0",x"ea",x"c2",x"50"),
  1076 => (x"1e",x"49",x"bf",x"97"),
  1077 => (x"d6",x"c1",x"49",x"c0"),
  1078 => (x"e9",x"c2",x"87",x"f5"),
  1079 => (x"78",x"de",x"48",x"f8"),
  1080 => (x"f4",x"d5",x"49",x"c1"),
  1081 => (x"fe",x"f6",x"26",x"87"),
  1082 => (x"4a",x"71",x"1e",x"87"),
  1083 => (x"c1",x"91",x"cb",x"49"),
  1084 => (x"c8",x"81",x"c5",x"dd"),
  1085 => (x"c2",x"48",x"11",x"81"),
  1086 => (x"c2",x"58",x"fc",x"e9"),
  1087 => (x"c0",x"48",x"fc",x"e9"),
  1088 => (x"d5",x"49",x"c1",x"78"),
  1089 => (x"4f",x"26",x"87",x"d3"),
  1090 => (x"c0",x"49",x"c0",x"1e"),
  1091 => (x"26",x"87",x"ca",x"fc"),
  1092 => (x"99",x"71",x"1e",x"4f"),
  1093 => (x"c1",x"87",x"d2",x"02"),
  1094 => (x"c0",x"48",x"da",x"de"),
  1095 => (x"c1",x"80",x"f7",x"50"),
  1096 => (x"c1",x"40",x"e9",x"c3"),
  1097 => (x"ce",x"78",x"fe",x"dc"),
  1098 => (x"d6",x"de",x"c1",x"87"),
  1099 => (x"f7",x"dc",x"c1",x"48"),
  1100 => (x"c1",x"80",x"fc",x"78"),
  1101 => (x"26",x"78",x"c8",x"c4"),
  1102 => (x"5b",x"5e",x"0e",x"4f"),
  1103 => (x"4c",x"71",x"0e",x"5c"),
  1104 => (x"c1",x"92",x"cb",x"4a"),
  1105 => (x"c8",x"82",x"c5",x"dd"),
  1106 => (x"a2",x"c9",x"49",x"a2"),
  1107 => (x"4b",x"6b",x"97",x"4b"),
  1108 => (x"49",x"69",x"97",x"1e"),
  1109 => (x"12",x"82",x"ca",x"1e"),
  1110 => (x"c5",x"e7",x"c0",x"49"),
  1111 => (x"d3",x"49",x"c0",x"87"),
  1112 => (x"49",x"74",x"87",x"f7"),
  1113 => (x"87",x"cc",x"f9",x"c0"),
  1114 => (x"f8",x"f4",x"8e",x"f8"),
  1115 => (x"1e",x"73",x"1e",x"87"),
  1116 => (x"ff",x"49",x"4b",x"71"),
  1117 => (x"49",x"73",x"87",x"c3"),
  1118 => (x"f4",x"87",x"fe",x"fe"),
  1119 => (x"73",x"1e",x"87",x"e9"),
  1120 => (x"c6",x"4b",x"71",x"1e"),
  1121 => (x"db",x"02",x"4a",x"a3"),
  1122 => (x"02",x"8a",x"c1",x"87"),
  1123 => (x"02",x"8a",x"87",x"d6"),
  1124 => (x"8a",x"87",x"da",x"c1"),
  1125 => (x"87",x"fc",x"c0",x"02"),
  1126 => (x"e1",x"c0",x"02",x"8a"),
  1127 => (x"cb",x"02",x"8a",x"87"),
  1128 => (x"87",x"db",x"c1",x"87"),
  1129 => (x"c0",x"fd",x"49",x"c7"),
  1130 => (x"87",x"de",x"c1",x"87"),
  1131 => (x"bf",x"fc",x"e9",x"c2"),
  1132 => (x"87",x"cb",x"c1",x"02"),
  1133 => (x"c2",x"88",x"c1",x"48"),
  1134 => (x"c1",x"58",x"c0",x"ea"),
  1135 => (x"ea",x"c2",x"87",x"c1"),
  1136 => (x"c0",x"02",x"bf",x"c0"),
  1137 => (x"e9",x"c2",x"87",x"f9"),
  1138 => (x"c1",x"48",x"bf",x"fc"),
  1139 => (x"c0",x"ea",x"c2",x"80"),
  1140 => (x"87",x"eb",x"c0",x"58"),
  1141 => (x"bf",x"fc",x"e9",x"c2"),
  1142 => (x"c2",x"89",x"c6",x"49"),
  1143 => (x"c0",x"59",x"c0",x"ea"),
  1144 => (x"da",x"03",x"a9",x"b7"),
  1145 => (x"fc",x"e9",x"c2",x"87"),
  1146 => (x"d2",x"78",x"c0",x"48"),
  1147 => (x"c0",x"ea",x"c2",x"87"),
  1148 => (x"87",x"cb",x"02",x"bf"),
  1149 => (x"bf",x"fc",x"e9",x"c2"),
  1150 => (x"c2",x"80",x"c6",x"48"),
  1151 => (x"c0",x"58",x"c0",x"ea"),
  1152 => (x"87",x"d5",x"d1",x"49"),
  1153 => (x"f6",x"c0",x"49",x"73"),
  1154 => (x"da",x"f2",x"87",x"ea"),
  1155 => (x"5b",x"5e",x"0e",x"87"),
  1156 => (x"4c",x"71",x"0e",x"5c"),
  1157 => (x"74",x"1e",x"66",x"cc"),
  1158 => (x"c1",x"93",x"cb",x"4b"),
  1159 => (x"c4",x"83",x"c5",x"dd"),
  1160 => (x"49",x"6a",x"4a",x"a3"),
  1161 => (x"87",x"d0",x"fa",x"fe"),
  1162 => (x"7b",x"e7",x"c2",x"c1"),
  1163 => (x"d4",x"49",x"a3",x"c8"),
  1164 => (x"a3",x"c9",x"51",x"66"),
  1165 => (x"51",x"66",x"d8",x"49"),
  1166 => (x"dc",x"49",x"a3",x"ca"),
  1167 => (x"f1",x"26",x"51",x"66"),
  1168 => (x"5e",x"0e",x"87",x"e3"),
  1169 => (x"0e",x"5d",x"5c",x"5b"),
  1170 => (x"d8",x"86",x"d0",x"ff"),
  1171 => (x"a6",x"c4",x"59",x"a6"),
  1172 => (x"c4",x"78",x"c0",x"48"),
  1173 => (x"66",x"c4",x"c1",x"80"),
  1174 => (x"c1",x"80",x"c4",x"78"),
  1175 => (x"c1",x"80",x"c4",x"78"),
  1176 => (x"c0",x"ea",x"c2",x"78"),
  1177 => (x"c2",x"78",x"c1",x"48"),
  1178 => (x"48",x"bf",x"f8",x"e9"),
  1179 => (x"cb",x"05",x"a8",x"de"),
  1180 => (x"87",x"e5",x"f3",x"87"),
  1181 => (x"a6",x"c8",x"49",x"70"),
  1182 => (x"87",x"e6",x"ce",x"59"),
  1183 => (x"e9",x"87",x"ed",x"e8"),
  1184 => (x"dc",x"e8",x"87",x"cf"),
  1185 => (x"c0",x"4c",x"70",x"87"),
  1186 => (x"c1",x"02",x"ac",x"fb"),
  1187 => (x"66",x"d4",x"87",x"d0"),
  1188 => (x"87",x"c2",x"c1",x"05"),
  1189 => (x"c1",x"1e",x"1e",x"c0"),
  1190 => (x"f8",x"de",x"c1",x"1e"),
  1191 => (x"fd",x"49",x"c0",x"1e"),
  1192 => (x"d0",x"c1",x"87",x"eb"),
  1193 => (x"82",x"c4",x"4a",x"66"),
  1194 => (x"81",x"c7",x"49",x"6a"),
  1195 => (x"1e",x"c1",x"51",x"74"),
  1196 => (x"49",x"6a",x"1e",x"d8"),
  1197 => (x"ec",x"e8",x"81",x"c8"),
  1198 => (x"c1",x"86",x"d8",x"87"),
  1199 => (x"c0",x"48",x"66",x"c4"),
  1200 => (x"87",x"c7",x"01",x"a8"),
  1201 => (x"c1",x"48",x"a6",x"c4"),
  1202 => (x"c1",x"87",x"ce",x"78"),
  1203 => (x"c1",x"48",x"66",x"c4"),
  1204 => (x"58",x"a6",x"cc",x"88"),
  1205 => (x"f8",x"e7",x"87",x"c3"),
  1206 => (x"48",x"a6",x"cc",x"87"),
  1207 => (x"9c",x"74",x"78",x"c2"),
  1208 => (x"87",x"fa",x"cc",x"02"),
  1209 => (x"c1",x"48",x"66",x"c4"),
  1210 => (x"03",x"a8",x"66",x"c8"),
  1211 => (x"d8",x"87",x"ef",x"cc"),
  1212 => (x"78",x"c0",x"48",x"a6"),
  1213 => (x"78",x"c0",x"80",x"c4"),
  1214 => (x"70",x"87",x"e6",x"e6"),
  1215 => (x"ac",x"d0",x"c1",x"4c"),
  1216 => (x"87",x"d7",x"c2",x"05"),
  1217 => (x"e9",x"7e",x"66",x"dc"),
  1218 => (x"49",x"70",x"87",x"ca"),
  1219 => (x"59",x"a6",x"e0",x"c0"),
  1220 => (x"70",x"87",x"ce",x"e6"),
  1221 => (x"ac",x"ec",x"c0",x"4c"),
  1222 => (x"87",x"ea",x"c1",x"05"),
  1223 => (x"cb",x"49",x"66",x"c4"),
  1224 => (x"66",x"c0",x"c1",x"91"),
  1225 => (x"4a",x"a1",x"c4",x"81"),
  1226 => (x"a1",x"c8",x"4d",x"6a"),
  1227 => (x"52",x"66",x"dc",x"4a"),
  1228 => (x"79",x"e9",x"c3",x"c1"),
  1229 => (x"70",x"87",x"ea",x"e5"),
  1230 => (x"d8",x"02",x"9c",x"4c"),
  1231 => (x"ac",x"fb",x"c0",x"87"),
  1232 => (x"74",x"87",x"d2",x"02"),
  1233 => (x"87",x"d9",x"e5",x"55"),
  1234 => (x"02",x"9c",x"4c",x"70"),
  1235 => (x"fb",x"c0",x"87",x"c7"),
  1236 => (x"ee",x"ff",x"05",x"ac"),
  1237 => (x"55",x"e0",x"c0",x"87"),
  1238 => (x"c0",x"55",x"c1",x"c2"),
  1239 => (x"66",x"d4",x"7d",x"97"),
  1240 => (x"05",x"a9",x"6e",x"49"),
  1241 => (x"66",x"c4",x"87",x"db"),
  1242 => (x"a8",x"66",x"c8",x"48"),
  1243 => (x"c4",x"87",x"ca",x"04"),
  1244 => (x"80",x"c1",x"48",x"66"),
  1245 => (x"c8",x"58",x"a6",x"c8"),
  1246 => (x"48",x"66",x"c8",x"87"),
  1247 => (x"a6",x"cc",x"88",x"c1"),
  1248 => (x"87",x"dd",x"e4",x"58"),
  1249 => (x"d0",x"c1",x"4c",x"70"),
  1250 => (x"87",x"c8",x"05",x"ac"),
  1251 => (x"c1",x"48",x"66",x"d0"),
  1252 => (x"58",x"a6",x"d4",x"80"),
  1253 => (x"02",x"ac",x"d0",x"c1"),
  1254 => (x"c0",x"87",x"e9",x"fd"),
  1255 => (x"d4",x"48",x"a6",x"e0"),
  1256 => (x"66",x"dc",x"78",x"66"),
  1257 => (x"66",x"e0",x"c0",x"48"),
  1258 => (x"c3",x"c9",x"05",x"a8"),
  1259 => (x"a6",x"e4",x"c0",x"87"),
  1260 => (x"7e",x"78",x"c0",x"48"),
  1261 => (x"fb",x"c0",x"48",x"74"),
  1262 => (x"a6",x"ec",x"c0",x"88"),
  1263 => (x"02",x"98",x"70",x"58"),
  1264 => (x"48",x"87",x"c8",x"c8"),
  1265 => (x"ec",x"c0",x"88",x"cb"),
  1266 => (x"98",x"70",x"58",x"a6"),
  1267 => (x"87",x"d0",x"c1",x"02"),
  1268 => (x"c0",x"88",x"c9",x"48"),
  1269 => (x"70",x"58",x"a6",x"ec"),
  1270 => (x"d6",x"c3",x"02",x"98"),
  1271 => (x"88",x"c4",x"48",x"87"),
  1272 => (x"58",x"a6",x"ec",x"c0"),
  1273 => (x"d0",x"02",x"98",x"70"),
  1274 => (x"88",x"c1",x"48",x"87"),
  1275 => (x"58",x"a6",x"ec",x"c0"),
  1276 => (x"c2",x"02",x"98",x"70"),
  1277 => (x"cc",x"c7",x"87",x"fd"),
  1278 => (x"48",x"a6",x"d8",x"87"),
  1279 => (x"e2",x"78",x"f0",x"c0"),
  1280 => (x"4c",x"70",x"87",x"df"),
  1281 => (x"02",x"ac",x"ec",x"c0"),
  1282 => (x"dc",x"87",x"c3",x"c0"),
  1283 => (x"ec",x"c0",x"5c",x"a6"),
  1284 => (x"87",x"cc",x"02",x"ac"),
  1285 => (x"70",x"87",x"ca",x"e2"),
  1286 => (x"ac",x"ec",x"c0",x"4c"),
  1287 => (x"87",x"f4",x"ff",x"05"),
  1288 => (x"02",x"ac",x"ec",x"c0"),
  1289 => (x"e1",x"87",x"c3",x"c0"),
  1290 => (x"66",x"d8",x"87",x"f7"),
  1291 => (x"49",x"66",x"d4",x"1e"),
  1292 => (x"49",x"66",x"d4",x"1e"),
  1293 => (x"f8",x"de",x"c1",x"1e"),
  1294 => (x"49",x"66",x"d4",x"1e"),
  1295 => (x"c0",x"87",x"ce",x"f7"),
  1296 => (x"dc",x"1e",x"ca",x"1e"),
  1297 => (x"91",x"cb",x"49",x"66"),
  1298 => (x"81",x"66",x"d8",x"c1"),
  1299 => (x"c4",x"48",x"a6",x"d8"),
  1300 => (x"66",x"d8",x"78",x"a1"),
  1301 => (x"cc",x"e2",x"49",x"bf"),
  1302 => (x"c0",x"86",x"d8",x"87"),
  1303 => (x"c1",x"06",x"a8",x"b7"),
  1304 => (x"1e",x"c1",x"87",x"c4"),
  1305 => (x"66",x"c8",x"1e",x"de"),
  1306 => (x"f8",x"e1",x"49",x"bf"),
  1307 => (x"70",x"86",x"c8",x"87"),
  1308 => (x"08",x"c0",x"48",x"49"),
  1309 => (x"58",x"a6",x"dc",x"88"),
  1310 => (x"06",x"a8",x"b7",x"c0"),
  1311 => (x"d8",x"87",x"e7",x"c0"),
  1312 => (x"b7",x"dd",x"48",x"66"),
  1313 => (x"87",x"de",x"03",x"a8"),
  1314 => (x"d8",x"49",x"bf",x"6e"),
  1315 => (x"e0",x"c0",x"81",x"66"),
  1316 => (x"49",x"66",x"d8",x"51"),
  1317 => (x"bf",x"6e",x"81",x"c1"),
  1318 => (x"51",x"c1",x"c2",x"81"),
  1319 => (x"c2",x"49",x"66",x"d8"),
  1320 => (x"81",x"bf",x"6e",x"81"),
  1321 => (x"66",x"cc",x"51",x"c0"),
  1322 => (x"d0",x"80",x"c1",x"48"),
  1323 => (x"7e",x"c1",x"58",x"a6"),
  1324 => (x"e2",x"87",x"d8",x"c4"),
  1325 => (x"a6",x"dc",x"87",x"de"),
  1326 => (x"87",x"d8",x"e2",x"58"),
  1327 => (x"58",x"a6",x"ec",x"c0"),
  1328 => (x"05",x"a8",x"ec",x"c0"),
  1329 => (x"c0",x"87",x"ca",x"c0"),
  1330 => (x"d8",x"48",x"a6",x"e8"),
  1331 => (x"c4",x"c0",x"78",x"66"),
  1332 => (x"cc",x"df",x"ff",x"87"),
  1333 => (x"49",x"66",x"c4",x"87"),
  1334 => (x"c0",x"c1",x"91",x"cb"),
  1335 => (x"80",x"71",x"48",x"66"),
  1336 => (x"4a",x"6e",x"7e",x"70"),
  1337 => (x"49",x"6e",x"82",x"c8"),
  1338 => (x"66",x"d8",x"81",x"ca"),
  1339 => (x"66",x"e8",x"c0",x"51"),
  1340 => (x"d8",x"81",x"c1",x"49"),
  1341 => (x"48",x"c1",x"89",x"66"),
  1342 => (x"49",x"70",x"30",x"71"),
  1343 => (x"97",x"71",x"89",x"c1"),
  1344 => (x"ed",x"ed",x"c2",x"7a"),
  1345 => (x"66",x"d8",x"49",x"bf"),
  1346 => (x"4a",x"6a",x"97",x"29"),
  1347 => (x"c0",x"98",x"71",x"48"),
  1348 => (x"6e",x"58",x"a6",x"f0"),
  1349 => (x"69",x"81",x"c4",x"49"),
  1350 => (x"66",x"e0",x"c0",x"4d"),
  1351 => (x"a8",x"66",x"dc",x"48"),
  1352 => (x"87",x"c8",x"c0",x"02"),
  1353 => (x"c0",x"48",x"a6",x"d8"),
  1354 => (x"87",x"c5",x"c0",x"78"),
  1355 => (x"c1",x"48",x"a6",x"d8"),
  1356 => (x"1e",x"66",x"d8",x"78"),
  1357 => (x"75",x"1e",x"e0",x"c0"),
  1358 => (x"e8",x"de",x"ff",x"49"),
  1359 => (x"70",x"86",x"c8",x"87"),
  1360 => (x"ac",x"b7",x"c0",x"4c"),
  1361 => (x"87",x"d4",x"c1",x"06"),
  1362 => (x"e0",x"c0",x"85",x"74"),
  1363 => (x"75",x"89",x"74",x"49"),
  1364 => (x"d6",x"d9",x"c1",x"4b"),
  1365 => (x"ed",x"fe",x"71",x"4a"),
  1366 => (x"85",x"c2",x"87",x"ce"),
  1367 => (x"48",x"66",x"e4",x"c0"),
  1368 => (x"e8",x"c0",x"80",x"c1"),
  1369 => (x"ec",x"c0",x"58",x"a6"),
  1370 => (x"81",x"c1",x"49",x"66"),
  1371 => (x"c0",x"02",x"a9",x"70"),
  1372 => (x"a6",x"d8",x"87",x"c8"),
  1373 => (x"c0",x"78",x"c0",x"48"),
  1374 => (x"a6",x"d8",x"87",x"c5"),
  1375 => (x"d8",x"78",x"c1",x"48"),
  1376 => (x"a4",x"c2",x"1e",x"66"),
  1377 => (x"48",x"e0",x"c0",x"49"),
  1378 => (x"49",x"70",x"88",x"71"),
  1379 => (x"ff",x"49",x"75",x"1e"),
  1380 => (x"c8",x"87",x"d2",x"dd"),
  1381 => (x"a8",x"b7",x"c0",x"86"),
  1382 => (x"87",x"c0",x"ff",x"01"),
  1383 => (x"02",x"66",x"e4",x"c0"),
  1384 => (x"6e",x"87",x"d1",x"c0"),
  1385 => (x"c0",x"81",x"c9",x"49"),
  1386 => (x"6e",x"51",x"66",x"e4"),
  1387 => (x"f9",x"c4",x"c1",x"48"),
  1388 => (x"87",x"cc",x"c0",x"78"),
  1389 => (x"81",x"c9",x"49",x"6e"),
  1390 => (x"48",x"6e",x"51",x"c2"),
  1391 => (x"78",x"ed",x"c5",x"c1"),
  1392 => (x"c6",x"c0",x"7e",x"c1"),
  1393 => (x"c8",x"dc",x"ff",x"87"),
  1394 => (x"6e",x"4c",x"70",x"87"),
  1395 => (x"87",x"f5",x"c0",x"02"),
  1396 => (x"c8",x"48",x"66",x"c4"),
  1397 => (x"c0",x"04",x"a8",x"66"),
  1398 => (x"66",x"c4",x"87",x"cb"),
  1399 => (x"c8",x"80",x"c1",x"48"),
  1400 => (x"e0",x"c0",x"58",x"a6"),
  1401 => (x"48",x"66",x"c8",x"87"),
  1402 => (x"a6",x"cc",x"88",x"c1"),
  1403 => (x"87",x"d5",x"c0",x"58"),
  1404 => (x"05",x"ac",x"c6",x"c1"),
  1405 => (x"cc",x"87",x"c8",x"c0"),
  1406 => (x"80",x"c1",x"48",x"66"),
  1407 => (x"ff",x"58",x"a6",x"d0"),
  1408 => (x"70",x"87",x"ce",x"db"),
  1409 => (x"48",x"66",x"d0",x"4c"),
  1410 => (x"a6",x"d4",x"80",x"c1"),
  1411 => (x"02",x"9c",x"74",x"58"),
  1412 => (x"c4",x"87",x"cb",x"c0"),
  1413 => (x"c8",x"c1",x"48",x"66"),
  1414 => (x"f3",x"04",x"a8",x"66"),
  1415 => (x"da",x"ff",x"87",x"d1"),
  1416 => (x"66",x"c4",x"87",x"e6"),
  1417 => (x"03",x"a8",x"c7",x"48"),
  1418 => (x"c2",x"87",x"e5",x"c0"),
  1419 => (x"c0",x"48",x"c0",x"ea"),
  1420 => (x"49",x"66",x"c4",x"78"),
  1421 => (x"c0",x"c1",x"91",x"cb"),
  1422 => (x"a1",x"c4",x"81",x"66"),
  1423 => (x"c0",x"4a",x"6a",x"4a"),
  1424 => (x"66",x"c4",x"79",x"52"),
  1425 => (x"c8",x"80",x"c1",x"48"),
  1426 => (x"a8",x"c7",x"58",x"a6"),
  1427 => (x"87",x"db",x"ff",x"04"),
  1428 => (x"e1",x"8e",x"d0",x"ff"),
  1429 => (x"20",x"3a",x"87",x"cd"),
  1430 => (x"1e",x"73",x"1e",x"00"),
  1431 => (x"02",x"9b",x"4b",x"71"),
  1432 => (x"e9",x"c2",x"87",x"c6"),
  1433 => (x"78",x"c0",x"48",x"fc"),
  1434 => (x"e9",x"c2",x"1e",x"c7"),
  1435 => (x"1e",x"49",x"bf",x"fc"),
  1436 => (x"1e",x"c5",x"dd",x"c1"),
  1437 => (x"bf",x"f8",x"e9",x"c2"),
  1438 => (x"87",x"c6",x"ef",x"49"),
  1439 => (x"e9",x"c2",x"86",x"cc"),
  1440 => (x"ea",x"49",x"bf",x"f8"),
  1441 => (x"9b",x"73",x"87",x"cb"),
  1442 => (x"c1",x"87",x"c8",x"02"),
  1443 => (x"c0",x"49",x"c5",x"dd"),
  1444 => (x"e0",x"87",x"f3",x"e5"),
  1445 => (x"c2",x"1e",x"87",x"d1"),
  1446 => (x"c0",x"48",x"cd",x"db"),
  1447 => (x"e8",x"de",x"c1",x"50"),
  1448 => (x"fb",x"c0",x"49",x"bf"),
  1449 => (x"48",x"c0",x"87",x"fc"),
  1450 => (x"c7",x"1e",x"4f",x"26"),
  1451 => (x"49",x"c1",x"87",x"e9"),
  1452 => (x"fe",x"87",x"e6",x"fe"),
  1453 => (x"70",x"87",x"c4",x"f0"),
  1454 => (x"87",x"cd",x"02",x"98"),
  1455 => (x"87",x"c1",x"f9",x"fe"),
  1456 => (x"c4",x"02",x"98",x"70"),
  1457 => (x"c2",x"4a",x"c1",x"87"),
  1458 => (x"72",x"4a",x"c0",x"87"),
  1459 => (x"87",x"ce",x"05",x"9a"),
  1460 => (x"db",x"c1",x"1e",x"c0"),
  1461 => (x"f1",x"c0",x"49",x"fe"),
  1462 => (x"86",x"c4",x"87",x"f0"),
  1463 => (x"c0",x"c1",x"87",x"fe"),
  1464 => (x"1e",x"c0",x"87",x"d5"),
  1465 => (x"49",x"c9",x"dc",x"c1"),
  1466 => (x"87",x"de",x"f1",x"c0"),
  1467 => (x"e5",x"fe",x"1e",x"c0"),
  1468 => (x"c0",x"49",x"70",x"87"),
  1469 => (x"c3",x"87",x"d3",x"f1"),
  1470 => (x"8e",x"f8",x"87",x"dc"),
  1471 => (x"44",x"53",x"4f",x"26"),
  1472 => (x"69",x"61",x"66",x"20"),
  1473 => (x"2e",x"64",x"65",x"6c"),
  1474 => (x"6f",x"6f",x"42",x"00"),
  1475 => (x"67",x"6e",x"69",x"74"),
  1476 => (x"00",x"2e",x"2e",x"2e"),
  1477 => (x"c9",x"e8",x"c0",x"1e"),
  1478 => (x"f4",x"f4",x"c0",x"87"),
  1479 => (x"26",x"87",x"f6",x"87"),
  1480 => (x"e9",x"c2",x"1e",x"4f"),
  1481 => (x"78",x"c0",x"48",x"fc"),
  1482 => (x"48",x"f8",x"e9",x"c2"),
  1483 => (x"f9",x"fd",x"78",x"c0"),
  1484 => (x"c0",x"87",x"e1",x"87"),
  1485 => (x"80",x"4f",x"26",x"48"),
  1486 => (x"69",x"78",x"45",x"20"),
  1487 => (x"20",x"80",x"00",x"74"),
  1488 => (x"6b",x"63",x"61",x"42"),
  1489 => (x"00",x"10",x"e9",x"00"),
  1490 => (x"00",x"2a",x"91",x"00"),
  1491 => (x"00",x"00",x"00",x"00"),
  1492 => (x"00",x"00",x"10",x"e9"),
  1493 => (x"00",x"00",x"2a",x"af"),
  1494 => (x"e9",x"00",x"00",x"00"),
  1495 => (x"cd",x"00",x"00",x"10"),
  1496 => (x"00",x"00",x"00",x"2a"),
  1497 => (x"10",x"e9",x"00",x"00"),
  1498 => (x"2a",x"eb",x"00",x"00"),
  1499 => (x"00",x"00",x"00",x"00"),
  1500 => (x"00",x"10",x"e9",x"00"),
  1501 => (x"00",x"2b",x"09",x"00"),
  1502 => (x"00",x"00",x"00",x"00"),
  1503 => (x"00",x"00",x"10",x"e9"),
  1504 => (x"00",x"00",x"2b",x"27"),
  1505 => (x"e9",x"00",x"00",x"00"),
  1506 => (x"45",x"00",x"00",x"10"),
  1507 => (x"00",x"00",x"00",x"2b"),
  1508 => (x"10",x"e9",x"00",x"00"),
  1509 => (x"00",x"00",x"00",x"00"),
  1510 => (x"00",x"00",x"00",x"00"),
  1511 => (x"00",x"11",x"7e",x"00"),
  1512 => (x"00",x"00",x"00",x"00"),
  1513 => (x"00",x"00",x"00",x"00"),
  1514 => (x"00",x"00",x"17",x"ac"),
  1515 => (x"54",x"4f",x"4f",x"42"),
  1516 => (x"20",x"20",x"20",x"20"),
  1517 => (x"00",x"4d",x"4f",x"52"),
  1518 => (x"64",x"61",x"6f",x"4c"),
  1519 => (x"00",x"2e",x"2a",x"20"),
  1520 => (x"48",x"f0",x"fe",x"1e"),
  1521 => (x"09",x"cd",x"78",x"c0"),
  1522 => (x"4f",x"26",x"09",x"79"),
  1523 => (x"f0",x"fe",x"1e",x"1e"),
  1524 => (x"26",x"48",x"7e",x"bf"),
  1525 => (x"fe",x"1e",x"4f",x"26"),
  1526 => (x"78",x"c1",x"48",x"f0"),
  1527 => (x"fe",x"1e",x"4f",x"26"),
  1528 => (x"78",x"c0",x"48",x"f0"),
  1529 => (x"71",x"1e",x"4f",x"26"),
  1530 => (x"52",x"52",x"c0",x"4a"),
  1531 => (x"5e",x"0e",x"4f",x"26"),
  1532 => (x"0e",x"5d",x"5c",x"5b"),
  1533 => (x"4d",x"71",x"86",x"f4"),
  1534 => (x"c1",x"7e",x"6d",x"97"),
  1535 => (x"6c",x"97",x"4c",x"a5"),
  1536 => (x"58",x"a6",x"c8",x"48"),
  1537 => (x"66",x"c4",x"48",x"6e"),
  1538 => (x"87",x"c5",x"05",x"a8"),
  1539 => (x"e6",x"c0",x"48",x"ff"),
  1540 => (x"87",x"ca",x"ff",x"87"),
  1541 => (x"97",x"49",x"a5",x"c2"),
  1542 => (x"a3",x"71",x"4b",x"6c"),
  1543 => (x"4b",x"6b",x"97",x"4b"),
  1544 => (x"6e",x"7e",x"6c",x"97"),
  1545 => (x"c8",x"80",x"c1",x"48"),
  1546 => (x"98",x"c7",x"58",x"a6"),
  1547 => (x"70",x"58",x"a6",x"cc"),
  1548 => (x"e1",x"fe",x"7c",x"97"),
  1549 => (x"f4",x"48",x"73",x"87"),
  1550 => (x"26",x"4d",x"26",x"8e"),
  1551 => (x"26",x"4b",x"26",x"4c"),
  1552 => (x"5b",x"5e",x"0e",x"4f"),
  1553 => (x"86",x"f4",x"0e",x"5c"),
  1554 => (x"66",x"d8",x"4c",x"71"),
  1555 => (x"9a",x"ff",x"c3",x"4a"),
  1556 => (x"97",x"4b",x"a4",x"c2"),
  1557 => (x"a1",x"73",x"49",x"6c"),
  1558 => (x"97",x"51",x"72",x"49"),
  1559 => (x"48",x"6e",x"7e",x"6c"),
  1560 => (x"a6",x"c8",x"80",x"c1"),
  1561 => (x"cc",x"98",x"c7",x"58"),
  1562 => (x"54",x"70",x"58",x"a6"),
  1563 => (x"ca",x"ff",x"8e",x"f4"),
  1564 => (x"fd",x"1e",x"1e",x"87"),
  1565 => (x"bf",x"e0",x"87",x"e8"),
  1566 => (x"e0",x"c0",x"49",x"4a"),
  1567 => (x"cb",x"02",x"99",x"c0"),
  1568 => (x"c2",x"1e",x"72",x"87"),
  1569 => (x"fe",x"49",x"e3",x"ed"),
  1570 => (x"86",x"c4",x"87",x"f7"),
  1571 => (x"70",x"87",x"fd",x"fc"),
  1572 => (x"87",x"c2",x"fd",x"7e"),
  1573 => (x"1e",x"4f",x"26",x"26"),
  1574 => (x"49",x"e3",x"ed",x"c2"),
  1575 => (x"c1",x"87",x"c7",x"fd"),
  1576 => (x"fc",x"49",x"f1",x"e1"),
  1577 => (x"d9",x"c5",x"87",x"da"),
  1578 => (x"0e",x"4f",x"26",x"87"),
  1579 => (x"5d",x"5c",x"5b",x"5e"),
  1580 => (x"c2",x"ee",x"c2",x"0e"),
  1581 => (x"e3",x"c1",x"4a",x"bf"),
  1582 => (x"4c",x"49",x"bf",x"ff"),
  1583 => (x"4d",x"71",x"bc",x"72"),
  1584 => (x"c0",x"87",x"db",x"fc"),
  1585 => (x"d0",x"49",x"74",x"4b"),
  1586 => (x"87",x"d5",x"02",x"99"),
  1587 => (x"99",x"d0",x"49",x"75"),
  1588 => (x"1e",x"c0",x"1e",x"71"),
  1589 => (x"4a",x"d1",x"ea",x"c1"),
  1590 => (x"49",x"12",x"82",x"73"),
  1591 => (x"c8",x"87",x"e4",x"c0"),
  1592 => (x"2d",x"2c",x"c1",x"86"),
  1593 => (x"04",x"ab",x"c8",x"83"),
  1594 => (x"fb",x"87",x"da",x"ff"),
  1595 => (x"e3",x"c1",x"87",x"e8"),
  1596 => (x"ee",x"c2",x"48",x"ff"),
  1597 => (x"26",x"78",x"bf",x"c2"),
  1598 => (x"26",x"4c",x"26",x"4d"),
  1599 => (x"00",x"4f",x"26",x"4b"),
  1600 => (x"1e",x"00",x"00",x"00"),
  1601 => (x"c8",x"48",x"d0",x"ff"),
  1602 => (x"d4",x"ff",x"78",x"e1"),
  1603 => (x"c4",x"78",x"c5",x"48"),
  1604 => (x"87",x"c3",x"02",x"66"),
  1605 => (x"c8",x"78",x"e0",x"c3"),
  1606 => (x"87",x"c6",x"02",x"66"),
  1607 => (x"c3",x"48",x"d4",x"ff"),
  1608 => (x"d4",x"ff",x"78",x"f0"),
  1609 => (x"ff",x"78",x"71",x"48"),
  1610 => (x"e1",x"c8",x"48",x"d0"),
  1611 => (x"78",x"e0",x"c0",x"78"),
  1612 => (x"5e",x"0e",x"4f",x"26"),
  1613 => (x"71",x"0e",x"5c",x"5b"),
  1614 => (x"e3",x"ed",x"c2",x"4c"),
  1615 => (x"87",x"ee",x"fa",x"49"),
  1616 => (x"b7",x"c0",x"4a",x"70"),
  1617 => (x"e3",x"c2",x"04",x"aa"),
  1618 => (x"aa",x"e0",x"c3",x"87"),
  1619 => (x"c1",x"87",x"c9",x"05"),
  1620 => (x"c1",x"48",x"f5",x"e7"),
  1621 => (x"87",x"d4",x"c2",x"78"),
  1622 => (x"05",x"aa",x"f0",x"c3"),
  1623 => (x"e7",x"c1",x"87",x"c9"),
  1624 => (x"78",x"c1",x"48",x"f1"),
  1625 => (x"c1",x"87",x"f5",x"c1"),
  1626 => (x"02",x"bf",x"f5",x"e7"),
  1627 => (x"4b",x"72",x"87",x"c7"),
  1628 => (x"c2",x"b3",x"c0",x"c2"),
  1629 => (x"74",x"4b",x"72",x"87"),
  1630 => (x"87",x"d1",x"05",x"9c"),
  1631 => (x"bf",x"f1",x"e7",x"c1"),
  1632 => (x"f5",x"e7",x"c1",x"1e"),
  1633 => (x"49",x"72",x"1e",x"bf"),
  1634 => (x"c8",x"87",x"f8",x"fd"),
  1635 => (x"f1",x"e7",x"c1",x"86"),
  1636 => (x"e0",x"c0",x"02",x"bf"),
  1637 => (x"c4",x"49",x"73",x"87"),
  1638 => (x"c1",x"91",x"29",x"b7"),
  1639 => (x"73",x"81",x"d1",x"e9"),
  1640 => (x"c2",x"9a",x"cf",x"4a"),
  1641 => (x"72",x"48",x"c1",x"92"),
  1642 => (x"ff",x"4a",x"70",x"30"),
  1643 => (x"69",x"48",x"72",x"ba"),
  1644 => (x"db",x"79",x"70",x"98"),
  1645 => (x"c4",x"49",x"73",x"87"),
  1646 => (x"c1",x"91",x"29",x"b7"),
  1647 => (x"73",x"81",x"d1",x"e9"),
  1648 => (x"c2",x"9a",x"cf",x"4a"),
  1649 => (x"72",x"48",x"c3",x"92"),
  1650 => (x"48",x"4a",x"70",x"30"),
  1651 => (x"79",x"70",x"b0",x"69"),
  1652 => (x"48",x"f5",x"e7",x"c1"),
  1653 => (x"e7",x"c1",x"78",x"c0"),
  1654 => (x"78",x"c0",x"48",x"f1"),
  1655 => (x"49",x"e3",x"ed",x"c2"),
  1656 => (x"70",x"87",x"cb",x"f8"),
  1657 => (x"aa",x"b7",x"c0",x"4a"),
  1658 => (x"87",x"dd",x"fd",x"03"),
  1659 => (x"c8",x"fc",x"48",x"c0"),
  1660 => (x"00",x"00",x"00",x"87"),
  1661 => (x"00",x"00",x"00",x"00"),
  1662 => (x"4a",x"71",x"1e",x"00"),
  1663 => (x"87",x"f2",x"fc",x"49"),
  1664 => (x"c0",x"1e",x"4f",x"26"),
  1665 => (x"c4",x"49",x"72",x"4a"),
  1666 => (x"d1",x"e9",x"c1",x"91"),
  1667 => (x"c1",x"79",x"c0",x"81"),
  1668 => (x"aa",x"b7",x"d0",x"82"),
  1669 => (x"26",x"87",x"ee",x"04"),
  1670 => (x"5b",x"5e",x"0e",x"4f"),
  1671 => (x"71",x"0e",x"5d",x"5c"),
  1672 => (x"87",x"fa",x"f6",x"4d"),
  1673 => (x"b7",x"c4",x"4a",x"75"),
  1674 => (x"e9",x"c1",x"92",x"2a"),
  1675 => (x"4c",x"75",x"82",x"d1"),
  1676 => (x"94",x"c2",x"9c",x"cf"),
  1677 => (x"74",x"4b",x"49",x"6a"),
  1678 => (x"c2",x"9b",x"c3",x"2b"),
  1679 => (x"70",x"30",x"74",x"48"),
  1680 => (x"74",x"bc",x"ff",x"4c"),
  1681 => (x"70",x"98",x"71",x"48"),
  1682 => (x"87",x"ca",x"f6",x"7a"),
  1683 => (x"e6",x"fa",x"48",x"73"),
  1684 => (x"00",x"00",x"00",x"87"),
  1685 => (x"00",x"00",x"00",x"00"),
  1686 => (x"00",x"00",x"00",x"00"),
  1687 => (x"00",x"00",x"00",x"00"),
  1688 => (x"00",x"00",x"00",x"00"),
  1689 => (x"00",x"00",x"00",x"00"),
  1690 => (x"00",x"00",x"00",x"00"),
  1691 => (x"00",x"00",x"00",x"00"),
  1692 => (x"00",x"00",x"00",x"00"),
  1693 => (x"00",x"00",x"00",x"00"),
  1694 => (x"00",x"00",x"00",x"00"),
  1695 => (x"00",x"00",x"00",x"00"),
  1696 => (x"00",x"00",x"00",x"00"),
  1697 => (x"00",x"00",x"00",x"00"),
  1698 => (x"00",x"00",x"00",x"00"),
  1699 => (x"00",x"00",x"00",x"00"),
  1700 => (x"26",x"1e",x"16",x"00"),
  1701 => (x"3d",x"36",x"2e",x"25"),
  1702 => (x"d0",x"ff",x"1e",x"3e"),
  1703 => (x"78",x"e1",x"c8",x"48"),
  1704 => (x"d4",x"ff",x"48",x"71"),
  1705 => (x"4f",x"26",x"78",x"08"),
  1706 => (x"48",x"d0",x"ff",x"1e"),
  1707 => (x"71",x"78",x"e1",x"c8"),
  1708 => (x"08",x"d4",x"ff",x"48"),
  1709 => (x"48",x"66",x"c4",x"78"),
  1710 => (x"78",x"08",x"d4",x"ff"),
  1711 => (x"71",x"1e",x"4f",x"26"),
  1712 => (x"49",x"66",x"c4",x"4a"),
  1713 => (x"ff",x"49",x"72",x"1e"),
  1714 => (x"d0",x"ff",x"87",x"de"),
  1715 => (x"78",x"e0",x"c0",x"48"),
  1716 => (x"1e",x"4f",x"26",x"26"),
  1717 => (x"66",x"c4",x"4a",x"71"),
  1718 => (x"a2",x"e0",x"c1",x"1e"),
  1719 => (x"87",x"c8",x"ff",x"49"),
  1720 => (x"c8",x"49",x"66",x"c8"),
  1721 => (x"d4",x"ff",x"29",x"b7"),
  1722 => (x"ff",x"78",x"71",x"48"),
  1723 => (x"e0",x"c0",x"48",x"d0"),
  1724 => (x"4f",x"26",x"26",x"78"),
  1725 => (x"4a",x"d4",x"ff",x"1e"),
  1726 => (x"ff",x"7a",x"ff",x"c3"),
  1727 => (x"e1",x"c8",x"48",x"d0"),
  1728 => (x"c2",x"7a",x"de",x"78"),
  1729 => (x"7a",x"bf",x"ed",x"ed"),
  1730 => (x"28",x"c8",x"48",x"49"),
  1731 => (x"48",x"71",x"7a",x"70"),
  1732 => (x"7a",x"70",x"28",x"d0"),
  1733 => (x"28",x"d8",x"48",x"71"),
  1734 => (x"d0",x"ff",x"7a",x"70"),
  1735 => (x"78",x"e0",x"c0",x"48"),
  1736 => (x"5e",x"0e",x"4f",x"26"),
  1737 => (x"0e",x"5d",x"5c",x"5b"),
  1738 => (x"ed",x"c2",x"4c",x"71"),
  1739 => (x"4b",x"4d",x"bf",x"ed"),
  1740 => (x"66",x"d0",x"2b",x"74"),
  1741 => (x"d4",x"83",x"c1",x"9b"),
  1742 => (x"c2",x"04",x"ab",x"66"),
  1743 => (x"74",x"4b",x"c0",x"87"),
  1744 => (x"49",x"66",x"d0",x"4a"),
  1745 => (x"b9",x"ff",x"31",x"72"),
  1746 => (x"48",x"73",x"99",x"75"),
  1747 => (x"4a",x"70",x"30",x"72"),
  1748 => (x"c2",x"b0",x"71",x"48"),
  1749 => (x"fe",x"58",x"f1",x"ed"),
  1750 => (x"4d",x"26",x"87",x"da"),
  1751 => (x"4b",x"26",x"4c",x"26"),
  1752 => (x"ff",x"1e",x"4f",x"26"),
  1753 => (x"c9",x"c8",x"48",x"d0"),
  1754 => (x"ff",x"48",x"71",x"78"),
  1755 => (x"26",x"78",x"08",x"d4"),
  1756 => (x"4a",x"71",x"1e",x"4f"),
  1757 => (x"ff",x"87",x"eb",x"49"),
  1758 => (x"78",x"c8",x"48",x"d0"),
  1759 => (x"73",x"1e",x"4f",x"26"),
  1760 => (x"c2",x"4b",x"71",x"1e"),
  1761 => (x"02",x"bf",x"fd",x"ed"),
  1762 => (x"eb",x"c2",x"87",x"c3"),
  1763 => (x"48",x"d0",x"ff",x"87"),
  1764 => (x"73",x"78",x"c9",x"c8"),
  1765 => (x"b1",x"e0",x"c0",x"49"),
  1766 => (x"71",x"48",x"d4",x"ff"),
  1767 => (x"f1",x"ed",x"c2",x"78"),
  1768 => (x"c8",x"78",x"c0",x"48"),
  1769 => (x"87",x"c5",x"02",x"66"),
  1770 => (x"c2",x"49",x"ff",x"c3"),
  1771 => (x"c2",x"49",x"c0",x"87"),
  1772 => (x"cc",x"59",x"f9",x"ed"),
  1773 => (x"87",x"c6",x"02",x"66"),
  1774 => (x"4a",x"d5",x"d5",x"c5"),
  1775 => (x"ff",x"cf",x"87",x"c4"),
  1776 => (x"ed",x"c2",x"4a",x"ff"),
  1777 => (x"ed",x"c2",x"5a",x"fd"),
  1778 => (x"78",x"c1",x"48",x"fd"),
  1779 => (x"4d",x"26",x"87",x"c4"),
  1780 => (x"4b",x"26",x"4c",x"26"),
  1781 => (x"5e",x"0e",x"4f",x"26"),
  1782 => (x"0e",x"5d",x"5c",x"5b"),
  1783 => (x"ed",x"c2",x"4a",x"71"),
  1784 => (x"72",x"4c",x"bf",x"f9"),
  1785 => (x"87",x"cb",x"02",x"9a"),
  1786 => (x"c1",x"91",x"c8",x"49"),
  1787 => (x"71",x"4b",x"f4",x"ed"),
  1788 => (x"c1",x"87",x"c4",x"83"),
  1789 => (x"c0",x"4b",x"f4",x"f1"),
  1790 => (x"74",x"49",x"13",x"4d"),
  1791 => (x"f5",x"ed",x"c2",x"99"),
  1792 => (x"d4",x"ff",x"b9",x"bf"),
  1793 => (x"c1",x"78",x"71",x"48"),
  1794 => (x"c8",x"85",x"2c",x"b7"),
  1795 => (x"e8",x"04",x"ad",x"b7"),
  1796 => (x"f1",x"ed",x"c2",x"87"),
  1797 => (x"80",x"c8",x"48",x"bf"),
  1798 => (x"58",x"f5",x"ed",x"c2"),
  1799 => (x"1e",x"87",x"ef",x"fe"),
  1800 => (x"4b",x"71",x"1e",x"73"),
  1801 => (x"02",x"9a",x"4a",x"13"),
  1802 => (x"49",x"72",x"87",x"cb"),
  1803 => (x"13",x"87",x"e7",x"fe"),
  1804 => (x"f5",x"05",x"9a",x"4a"),
  1805 => (x"87",x"da",x"fe",x"87"),
  1806 => (x"f1",x"ed",x"c2",x"1e"),
  1807 => (x"ed",x"c2",x"49",x"bf"),
  1808 => (x"a1",x"c1",x"48",x"f1"),
  1809 => (x"b7",x"c0",x"c4",x"78"),
  1810 => (x"87",x"db",x"03",x"a9"),
  1811 => (x"c2",x"48",x"d4",x"ff"),
  1812 => (x"78",x"bf",x"f5",x"ed"),
  1813 => (x"bf",x"f1",x"ed",x"c2"),
  1814 => (x"f1",x"ed",x"c2",x"49"),
  1815 => (x"78",x"a1",x"c1",x"48"),
  1816 => (x"a9",x"b7",x"c0",x"c4"),
  1817 => (x"ff",x"87",x"e5",x"04"),
  1818 => (x"78",x"c8",x"48",x"d0"),
  1819 => (x"48",x"fd",x"ed",x"c2"),
  1820 => (x"4f",x"26",x"78",x"c0"),
  1821 => (x"00",x"00",x"00",x"00"),
  1822 => (x"00",x"00",x"00",x"00"),
  1823 => (x"5f",x"00",x"00",x"00"),
  1824 => (x"00",x"00",x"00",x"5f"),
  1825 => (x"00",x"03",x"03",x"00"),
  1826 => (x"00",x"00",x"03",x"03"),
  1827 => (x"14",x"7f",x"7f",x"14"),
  1828 => (x"00",x"14",x"7f",x"7f"),
  1829 => (x"6b",x"2e",x"24",x"00"),
  1830 => (x"00",x"12",x"3a",x"6b"),
  1831 => (x"18",x"36",x"6a",x"4c"),
  1832 => (x"00",x"32",x"56",x"6c"),
  1833 => (x"59",x"4f",x"7e",x"30"),
  1834 => (x"40",x"68",x"3a",x"77"),
  1835 => (x"07",x"04",x"00",x"00"),
  1836 => (x"00",x"00",x"00",x"03"),
  1837 => (x"3e",x"1c",x"00",x"00"),
  1838 => (x"00",x"00",x"41",x"63"),
  1839 => (x"63",x"41",x"00",x"00"),
  1840 => (x"00",x"00",x"1c",x"3e"),
  1841 => (x"1c",x"3e",x"2a",x"08"),
  1842 => (x"08",x"2a",x"3e",x"1c"),
  1843 => (x"3e",x"08",x"08",x"00"),
  1844 => (x"00",x"08",x"08",x"3e"),
  1845 => (x"e0",x"80",x"00",x"00"),
  1846 => (x"00",x"00",x"00",x"60"),
  1847 => (x"08",x"08",x"08",x"00"),
  1848 => (x"00",x"08",x"08",x"08"),
  1849 => (x"60",x"00",x"00",x"00"),
  1850 => (x"00",x"00",x"00",x"60"),
  1851 => (x"18",x"30",x"60",x"40"),
  1852 => (x"01",x"03",x"06",x"0c"),
  1853 => (x"59",x"7f",x"3e",x"00"),
  1854 => (x"00",x"3e",x"7f",x"4d"),
  1855 => (x"7f",x"06",x"04",x"00"),
  1856 => (x"00",x"00",x"00",x"7f"),
  1857 => (x"71",x"63",x"42",x"00"),
  1858 => (x"00",x"46",x"4f",x"59"),
  1859 => (x"49",x"63",x"22",x"00"),
  1860 => (x"00",x"36",x"7f",x"49"),
  1861 => (x"13",x"16",x"1c",x"18"),
  1862 => (x"00",x"10",x"7f",x"7f"),
  1863 => (x"45",x"67",x"27",x"00"),
  1864 => (x"00",x"39",x"7d",x"45"),
  1865 => (x"4b",x"7e",x"3c",x"00"),
  1866 => (x"00",x"30",x"79",x"49"),
  1867 => (x"71",x"01",x"01",x"00"),
  1868 => (x"00",x"07",x"0f",x"79"),
  1869 => (x"49",x"7f",x"36",x"00"),
  1870 => (x"00",x"36",x"7f",x"49"),
  1871 => (x"49",x"4f",x"06",x"00"),
  1872 => (x"00",x"1e",x"3f",x"69"),
  1873 => (x"66",x"00",x"00",x"00"),
  1874 => (x"00",x"00",x"00",x"66"),
  1875 => (x"e6",x"80",x"00",x"00"),
  1876 => (x"00",x"00",x"00",x"66"),
  1877 => (x"14",x"08",x"08",x"00"),
  1878 => (x"00",x"22",x"22",x"14"),
  1879 => (x"14",x"14",x"14",x"00"),
  1880 => (x"00",x"14",x"14",x"14"),
  1881 => (x"14",x"22",x"22",x"00"),
  1882 => (x"00",x"08",x"08",x"14"),
  1883 => (x"51",x"03",x"02",x"00"),
  1884 => (x"00",x"06",x"0f",x"59"),
  1885 => (x"5d",x"41",x"7f",x"3e"),
  1886 => (x"00",x"1e",x"1f",x"55"),
  1887 => (x"09",x"7f",x"7e",x"00"),
  1888 => (x"00",x"7e",x"7f",x"09"),
  1889 => (x"49",x"7f",x"7f",x"00"),
  1890 => (x"00",x"36",x"7f",x"49"),
  1891 => (x"63",x"3e",x"1c",x"00"),
  1892 => (x"00",x"41",x"41",x"41"),
  1893 => (x"41",x"7f",x"7f",x"00"),
  1894 => (x"00",x"1c",x"3e",x"63"),
  1895 => (x"49",x"7f",x"7f",x"00"),
  1896 => (x"00",x"41",x"41",x"49"),
  1897 => (x"09",x"7f",x"7f",x"00"),
  1898 => (x"00",x"01",x"01",x"09"),
  1899 => (x"41",x"7f",x"3e",x"00"),
  1900 => (x"00",x"7a",x"7b",x"49"),
  1901 => (x"08",x"7f",x"7f",x"00"),
  1902 => (x"00",x"7f",x"7f",x"08"),
  1903 => (x"7f",x"41",x"00",x"00"),
  1904 => (x"00",x"00",x"41",x"7f"),
  1905 => (x"40",x"60",x"20",x"00"),
  1906 => (x"00",x"3f",x"7f",x"40"),
  1907 => (x"1c",x"08",x"7f",x"7f"),
  1908 => (x"00",x"41",x"63",x"36"),
  1909 => (x"40",x"7f",x"7f",x"00"),
  1910 => (x"00",x"40",x"40",x"40"),
  1911 => (x"0c",x"06",x"7f",x"7f"),
  1912 => (x"00",x"7f",x"7f",x"06"),
  1913 => (x"0c",x"06",x"7f",x"7f"),
  1914 => (x"00",x"7f",x"7f",x"18"),
  1915 => (x"41",x"7f",x"3e",x"00"),
  1916 => (x"00",x"3e",x"7f",x"41"),
  1917 => (x"09",x"7f",x"7f",x"00"),
  1918 => (x"00",x"06",x"0f",x"09"),
  1919 => (x"61",x"41",x"7f",x"3e"),
  1920 => (x"00",x"40",x"7e",x"7f"),
  1921 => (x"09",x"7f",x"7f",x"00"),
  1922 => (x"00",x"66",x"7f",x"19"),
  1923 => (x"4d",x"6f",x"26",x"00"),
  1924 => (x"00",x"32",x"7b",x"59"),
  1925 => (x"7f",x"01",x"01",x"00"),
  1926 => (x"00",x"01",x"01",x"7f"),
  1927 => (x"40",x"7f",x"3f",x"00"),
  1928 => (x"00",x"3f",x"7f",x"40"),
  1929 => (x"70",x"3f",x"0f",x"00"),
  1930 => (x"00",x"0f",x"3f",x"70"),
  1931 => (x"18",x"30",x"7f",x"7f"),
  1932 => (x"00",x"7f",x"7f",x"30"),
  1933 => (x"1c",x"36",x"63",x"41"),
  1934 => (x"41",x"63",x"36",x"1c"),
  1935 => (x"7c",x"06",x"03",x"01"),
  1936 => (x"01",x"03",x"06",x"7c"),
  1937 => (x"4d",x"59",x"71",x"61"),
  1938 => (x"00",x"41",x"43",x"47"),
  1939 => (x"7f",x"7f",x"00",x"00"),
  1940 => (x"00",x"00",x"41",x"41"),
  1941 => (x"0c",x"06",x"03",x"01"),
  1942 => (x"40",x"60",x"30",x"18"),
  1943 => (x"41",x"41",x"00",x"00"),
  1944 => (x"00",x"00",x"7f",x"7f"),
  1945 => (x"03",x"06",x"0c",x"08"),
  1946 => (x"00",x"08",x"0c",x"06"),
  1947 => (x"80",x"80",x"80",x"80"),
  1948 => (x"00",x"80",x"80",x"80"),
  1949 => (x"03",x"00",x"00",x"00"),
  1950 => (x"00",x"00",x"04",x"07"),
  1951 => (x"54",x"74",x"20",x"00"),
  1952 => (x"00",x"78",x"7c",x"54"),
  1953 => (x"44",x"7f",x"7f",x"00"),
  1954 => (x"00",x"38",x"7c",x"44"),
  1955 => (x"44",x"7c",x"38",x"00"),
  1956 => (x"00",x"00",x"44",x"44"),
  1957 => (x"44",x"7c",x"38",x"00"),
  1958 => (x"00",x"7f",x"7f",x"44"),
  1959 => (x"54",x"7c",x"38",x"00"),
  1960 => (x"00",x"18",x"5c",x"54"),
  1961 => (x"7f",x"7e",x"04",x"00"),
  1962 => (x"00",x"00",x"05",x"05"),
  1963 => (x"a4",x"bc",x"18",x"00"),
  1964 => (x"00",x"7c",x"fc",x"a4"),
  1965 => (x"04",x"7f",x"7f",x"00"),
  1966 => (x"00",x"78",x"7c",x"04"),
  1967 => (x"3d",x"00",x"00",x"00"),
  1968 => (x"00",x"00",x"40",x"7d"),
  1969 => (x"80",x"80",x"80",x"00"),
  1970 => (x"00",x"00",x"7d",x"fd"),
  1971 => (x"10",x"7f",x"7f",x"00"),
  1972 => (x"00",x"44",x"6c",x"38"),
  1973 => (x"3f",x"00",x"00",x"00"),
  1974 => (x"00",x"00",x"40",x"7f"),
  1975 => (x"18",x"0c",x"7c",x"7c"),
  1976 => (x"00",x"78",x"7c",x"0c"),
  1977 => (x"04",x"7c",x"7c",x"00"),
  1978 => (x"00",x"78",x"7c",x"04"),
  1979 => (x"44",x"7c",x"38",x"00"),
  1980 => (x"00",x"38",x"7c",x"44"),
  1981 => (x"24",x"fc",x"fc",x"00"),
  1982 => (x"00",x"18",x"3c",x"24"),
  1983 => (x"24",x"3c",x"18",x"00"),
  1984 => (x"00",x"fc",x"fc",x"24"),
  1985 => (x"04",x"7c",x"7c",x"00"),
  1986 => (x"00",x"08",x"0c",x"04"),
  1987 => (x"54",x"5c",x"48",x"00"),
  1988 => (x"00",x"20",x"74",x"54"),
  1989 => (x"7f",x"3f",x"04",x"00"),
  1990 => (x"00",x"00",x"44",x"44"),
  1991 => (x"40",x"7c",x"3c",x"00"),
  1992 => (x"00",x"7c",x"7c",x"40"),
  1993 => (x"60",x"3c",x"1c",x"00"),
  1994 => (x"00",x"1c",x"3c",x"60"),
  1995 => (x"30",x"60",x"7c",x"3c"),
  1996 => (x"00",x"3c",x"7c",x"60"),
  1997 => (x"10",x"38",x"6c",x"44"),
  1998 => (x"00",x"44",x"6c",x"38"),
  1999 => (x"e0",x"bc",x"1c",x"00"),
  2000 => (x"00",x"1c",x"3c",x"60"),
  2001 => (x"74",x"64",x"44",x"00"),
  2002 => (x"00",x"44",x"4c",x"5c"),
  2003 => (x"3e",x"08",x"08",x"00"),
  2004 => (x"00",x"41",x"41",x"77"),
  2005 => (x"7f",x"00",x"00",x"00"),
  2006 => (x"00",x"00",x"00",x"7f"),
  2007 => (x"77",x"41",x"41",x"00"),
  2008 => (x"00",x"08",x"08",x"3e"),
  2009 => (x"03",x"01",x"01",x"02"),
  2010 => (x"00",x"01",x"02",x"02"),
  2011 => (x"7f",x"7f",x"7f",x"7f"),
  2012 => (x"00",x"7f",x"7f",x"7f"),
  2013 => (x"1c",x"1c",x"08",x"08"),
  2014 => (x"7f",x"7f",x"3e",x"3e"),
  2015 => (x"3e",x"3e",x"7f",x"7f"),
  2016 => (x"08",x"08",x"1c",x"1c"),
  2017 => (x"7c",x"18",x"10",x"00"),
  2018 => (x"00",x"10",x"18",x"7c"),
  2019 => (x"7c",x"30",x"10",x"00"),
  2020 => (x"00",x"10",x"30",x"7c"),
  2021 => (x"60",x"60",x"30",x"10"),
  2022 => (x"00",x"06",x"1e",x"78"),
  2023 => (x"18",x"3c",x"66",x"42"),
  2024 => (x"00",x"42",x"66",x"3c"),
  2025 => (x"c2",x"6a",x"38",x"78"),
  2026 => (x"00",x"38",x"6c",x"c6"),
  2027 => (x"60",x"00",x"00",x"60"),
  2028 => (x"00",x"60",x"00",x"00"),
  2029 => (x"5c",x"5b",x"5e",x"0e"),
  2030 => (x"71",x"1e",x"0e",x"5d"),
  2031 => (x"ce",x"ee",x"c2",x"4c"),
  2032 => (x"4b",x"c0",x"4d",x"bf"),
  2033 => (x"ab",x"74",x"1e",x"c0"),
  2034 => (x"c4",x"87",x"c7",x"02"),
  2035 => (x"78",x"c0",x"48",x"a6"),
  2036 => (x"a6",x"c4",x"87",x"c5"),
  2037 => (x"c4",x"78",x"c1",x"48"),
  2038 => (x"49",x"73",x"1e",x"66"),
  2039 => (x"c8",x"87",x"df",x"ee"),
  2040 => (x"49",x"e0",x"c0",x"86"),
  2041 => (x"c4",x"87",x"ef",x"ef"),
  2042 => (x"49",x"6a",x"4a",x"a5"),
  2043 => (x"f1",x"87",x"f0",x"f0"),
  2044 => (x"85",x"cb",x"87",x"c6"),
  2045 => (x"b7",x"c8",x"83",x"c1"),
  2046 => (x"c7",x"ff",x"04",x"ab"),
  2047 => (x"4d",x"26",x"26",x"87"),
  2048 => (x"4b",x"26",x"4c",x"26"),
  2049 => (x"71",x"1e",x"4f",x"26"),
  2050 => (x"d2",x"ee",x"c2",x"4a"),
  2051 => (x"d2",x"ee",x"c2",x"5a"),
  2052 => (x"49",x"78",x"c7",x"48"),
  2053 => (x"26",x"87",x"dd",x"fe"),
  2054 => (x"1e",x"73",x"1e",x"4f"),
  2055 => (x"b7",x"c0",x"4a",x"71"),
  2056 => (x"87",x"d3",x"03",x"aa"),
  2057 => (x"bf",x"f0",x"ce",x"c2"),
  2058 => (x"c1",x"87",x"c4",x"05"),
  2059 => (x"c0",x"87",x"c2",x"4b"),
  2060 => (x"f4",x"ce",x"c2",x"4b"),
  2061 => (x"c2",x"87",x"c4",x"5b"),
  2062 => (x"c2",x"5a",x"f4",x"ce"),
  2063 => (x"4a",x"bf",x"f0",x"ce"),
  2064 => (x"c0",x"c1",x"9a",x"c1"),
  2065 => (x"e8",x"ec",x"49",x"a2"),
  2066 => (x"c2",x"48",x"fc",x"87"),
  2067 => (x"78",x"bf",x"f0",x"ce"),
  2068 => (x"1e",x"87",x"ef",x"fe"),
  2069 => (x"66",x"c4",x"4a",x"71"),
  2070 => (x"e9",x"49",x"72",x"1e"),
  2071 => (x"26",x"26",x"87",x"f5"),
  2072 => (x"ce",x"c2",x"1e",x"4f"),
  2073 => (x"e6",x"49",x"bf",x"f0"),
  2074 => (x"ee",x"c2",x"87",x"cf"),
  2075 => (x"bf",x"e8",x"48",x"c6"),
  2076 => (x"c2",x"ee",x"c2",x"78"),
  2077 => (x"78",x"bf",x"ec",x"48"),
  2078 => (x"bf",x"c6",x"ee",x"c2"),
  2079 => (x"ff",x"c3",x"49",x"4a"),
  2080 => (x"2a",x"b7",x"c8",x"99"),
  2081 => (x"b0",x"71",x"48",x"72"),
  2082 => (x"58",x"ce",x"ee",x"c2"),
  2083 => (x"5e",x"0e",x"4f",x"26"),
  2084 => (x"0e",x"5d",x"5c",x"5b"),
  2085 => (x"c8",x"ff",x"4b",x"71"),
  2086 => (x"c1",x"ee",x"c2",x"87"),
  2087 => (x"73",x"50",x"c0",x"48"),
  2088 => (x"87",x"f5",x"e5",x"49"),
  2089 => (x"c2",x"4c",x"49",x"70"),
  2090 => (x"49",x"ee",x"cb",x"9c"),
  2091 => (x"70",x"87",x"c9",x"cc"),
  2092 => (x"ee",x"c2",x"4d",x"49"),
  2093 => (x"05",x"bf",x"97",x"c1"),
  2094 => (x"d0",x"87",x"e2",x"c1"),
  2095 => (x"ee",x"c2",x"49",x"66"),
  2096 => (x"05",x"99",x"bf",x"ca"),
  2097 => (x"66",x"d4",x"87",x"d6"),
  2098 => (x"c2",x"ee",x"c2",x"49"),
  2099 => (x"cb",x"05",x"99",x"bf"),
  2100 => (x"e5",x"49",x"73",x"87"),
  2101 => (x"98",x"70",x"87",x"c3"),
  2102 => (x"87",x"c1",x"c1",x"02"),
  2103 => (x"c0",x"fe",x"4c",x"c1"),
  2104 => (x"cb",x"49",x"75",x"87"),
  2105 => (x"98",x"70",x"87",x"de"),
  2106 => (x"c2",x"87",x"c6",x"02"),
  2107 => (x"c1",x"48",x"c1",x"ee"),
  2108 => (x"c1",x"ee",x"c2",x"50"),
  2109 => (x"c0",x"05",x"bf",x"97"),
  2110 => (x"ee",x"c2",x"87",x"e3"),
  2111 => (x"d0",x"49",x"bf",x"ca"),
  2112 => (x"ff",x"05",x"99",x"66"),
  2113 => (x"ee",x"c2",x"87",x"d6"),
  2114 => (x"d4",x"49",x"bf",x"c2"),
  2115 => (x"ff",x"05",x"99",x"66"),
  2116 => (x"49",x"73",x"87",x"ca"),
  2117 => (x"70",x"87",x"c2",x"e4"),
  2118 => (x"ff",x"fe",x"05",x"98"),
  2119 => (x"fb",x"48",x"74",x"87"),
  2120 => (x"5e",x"0e",x"87",x"dc"),
  2121 => (x"0e",x"5d",x"5c",x"5b"),
  2122 => (x"4d",x"c0",x"86",x"f4"),
  2123 => (x"7e",x"bf",x"ec",x"4c"),
  2124 => (x"c2",x"48",x"a6",x"c4"),
  2125 => (x"78",x"bf",x"ce",x"ee"),
  2126 => (x"1e",x"c0",x"1e",x"c1"),
  2127 => (x"cd",x"fd",x"49",x"c7"),
  2128 => (x"70",x"86",x"c8",x"87"),
  2129 => (x"87",x"cd",x"02",x"98"),
  2130 => (x"cc",x"fb",x"49",x"ff"),
  2131 => (x"49",x"da",x"c1",x"87"),
  2132 => (x"c1",x"87",x"c6",x"e3"),
  2133 => (x"c1",x"ee",x"c2",x"4d"),
  2134 => (x"c3",x"02",x"bf",x"97"),
  2135 => (x"87",x"ee",x"d5",x"87"),
  2136 => (x"bf",x"c6",x"ee",x"c2"),
  2137 => (x"f0",x"ce",x"c2",x"4b"),
  2138 => (x"d9",x"c1",x"05",x"bf"),
  2139 => (x"48",x"a6",x"c4",x"87"),
  2140 => (x"78",x"c0",x"c0",x"c8"),
  2141 => (x"7e",x"dc",x"ce",x"c2"),
  2142 => (x"49",x"bf",x"97",x"6e"),
  2143 => (x"80",x"c1",x"48",x"6e"),
  2144 => (x"e2",x"71",x"7e",x"70"),
  2145 => (x"98",x"70",x"87",x"d3"),
  2146 => (x"c4",x"87",x"c3",x"02"),
  2147 => (x"66",x"c4",x"b3",x"66"),
  2148 => (x"28",x"b7",x"c1",x"48"),
  2149 => (x"70",x"58",x"a6",x"c8"),
  2150 => (x"db",x"ff",x"05",x"98"),
  2151 => (x"49",x"fd",x"c3",x"87"),
  2152 => (x"c3",x"87",x"f6",x"e1"),
  2153 => (x"f0",x"e1",x"49",x"fa"),
  2154 => (x"c3",x"49",x"73",x"87"),
  2155 => (x"1e",x"71",x"99",x"ff"),
  2156 => (x"de",x"fa",x"49",x"c0"),
  2157 => (x"c8",x"49",x"73",x"87"),
  2158 => (x"1e",x"71",x"29",x"b7"),
  2159 => (x"d2",x"fa",x"49",x"c1"),
  2160 => (x"c5",x"86",x"c8",x"87"),
  2161 => (x"ee",x"c2",x"87",x"ff"),
  2162 => (x"9b",x"4b",x"bf",x"ca"),
  2163 => (x"c2",x"87",x"dd",x"02"),
  2164 => (x"49",x"bf",x"ec",x"ce"),
  2165 => (x"70",x"87",x"ed",x"c7"),
  2166 => (x"87",x"c4",x"05",x"98"),
  2167 => (x"87",x"d2",x"4b",x"c0"),
  2168 => (x"c7",x"49",x"e0",x"c2"),
  2169 => (x"ce",x"c2",x"87",x"d2"),
  2170 => (x"87",x"c6",x"58",x"f0"),
  2171 => (x"48",x"ec",x"ce",x"c2"),
  2172 => (x"49",x"73",x"78",x"c0"),
  2173 => (x"cd",x"05",x"99",x"c2"),
  2174 => (x"49",x"eb",x"c3",x"87"),
  2175 => (x"70",x"87",x"da",x"e0"),
  2176 => (x"02",x"99",x"c2",x"49"),
  2177 => (x"4c",x"fb",x"87",x"c2"),
  2178 => (x"99",x"c1",x"49",x"73"),
  2179 => (x"c3",x"87",x"cd",x"05"),
  2180 => (x"c4",x"e0",x"49",x"f4"),
  2181 => (x"c2",x"49",x"70",x"87"),
  2182 => (x"87",x"c2",x"02",x"99"),
  2183 => (x"49",x"73",x"4c",x"fa"),
  2184 => (x"ce",x"05",x"99",x"c8"),
  2185 => (x"49",x"f5",x"c3",x"87"),
  2186 => (x"87",x"ed",x"df",x"ff"),
  2187 => (x"99",x"c2",x"49",x"70"),
  2188 => (x"c2",x"87",x"d5",x"02"),
  2189 => (x"02",x"bf",x"d2",x"ee"),
  2190 => (x"c1",x"48",x"87",x"ca"),
  2191 => (x"d6",x"ee",x"c2",x"88"),
  2192 => (x"87",x"c2",x"c0",x"58"),
  2193 => (x"4d",x"c1",x"4c",x"ff"),
  2194 => (x"99",x"c4",x"49",x"73"),
  2195 => (x"c3",x"87",x"ce",x"05"),
  2196 => (x"df",x"ff",x"49",x"f2"),
  2197 => (x"49",x"70",x"87",x"c3"),
  2198 => (x"dc",x"02",x"99",x"c2"),
  2199 => (x"d2",x"ee",x"c2",x"87"),
  2200 => (x"c7",x"48",x"7e",x"bf"),
  2201 => (x"c0",x"03",x"a8",x"b7"),
  2202 => (x"48",x"6e",x"87",x"cb"),
  2203 => (x"ee",x"c2",x"80",x"c1"),
  2204 => (x"c2",x"c0",x"58",x"d6"),
  2205 => (x"c1",x"4c",x"fe",x"87"),
  2206 => (x"49",x"fd",x"c3",x"4d"),
  2207 => (x"87",x"d9",x"de",x"ff"),
  2208 => (x"99",x"c2",x"49",x"70"),
  2209 => (x"87",x"d5",x"c0",x"02"),
  2210 => (x"bf",x"d2",x"ee",x"c2"),
  2211 => (x"87",x"c9",x"c0",x"02"),
  2212 => (x"48",x"d2",x"ee",x"c2"),
  2213 => (x"c2",x"c0",x"78",x"c0"),
  2214 => (x"c1",x"4c",x"fd",x"87"),
  2215 => (x"49",x"fa",x"c3",x"4d"),
  2216 => (x"87",x"f5",x"dd",x"ff"),
  2217 => (x"99",x"c2",x"49",x"70"),
  2218 => (x"87",x"d9",x"c0",x"02"),
  2219 => (x"bf",x"d2",x"ee",x"c2"),
  2220 => (x"a8",x"b7",x"c7",x"48"),
  2221 => (x"87",x"c9",x"c0",x"03"),
  2222 => (x"48",x"d2",x"ee",x"c2"),
  2223 => (x"c2",x"c0",x"78",x"c7"),
  2224 => (x"c1",x"4c",x"fc",x"87"),
  2225 => (x"ac",x"b7",x"c0",x"4d"),
  2226 => (x"87",x"d1",x"c0",x"03"),
  2227 => (x"c1",x"4a",x"66",x"c4"),
  2228 => (x"02",x"6a",x"82",x"d8"),
  2229 => (x"6a",x"87",x"c6",x"c0"),
  2230 => (x"73",x"49",x"74",x"4b"),
  2231 => (x"c3",x"1e",x"c0",x"0f"),
  2232 => (x"da",x"c1",x"1e",x"f0"),
  2233 => (x"87",x"e6",x"f6",x"49"),
  2234 => (x"98",x"70",x"86",x"c8"),
  2235 => (x"87",x"e2",x"c0",x"02"),
  2236 => (x"c2",x"48",x"a6",x"c8"),
  2237 => (x"78",x"bf",x"d2",x"ee"),
  2238 => (x"cb",x"49",x"66",x"c8"),
  2239 => (x"48",x"66",x"c4",x"91"),
  2240 => (x"7e",x"70",x"80",x"71"),
  2241 => (x"c0",x"02",x"bf",x"6e"),
  2242 => (x"bf",x"6e",x"87",x"c8"),
  2243 => (x"49",x"66",x"c8",x"4b"),
  2244 => (x"9d",x"75",x"0f",x"73"),
  2245 => (x"87",x"c8",x"c0",x"02"),
  2246 => (x"bf",x"d2",x"ee",x"c2"),
  2247 => (x"87",x"d4",x"f2",x"49"),
  2248 => (x"bf",x"f4",x"ce",x"c2"),
  2249 => (x"87",x"dd",x"c0",x"02"),
  2250 => (x"87",x"d8",x"c2",x"49"),
  2251 => (x"c0",x"02",x"98",x"70"),
  2252 => (x"ee",x"c2",x"87",x"d3"),
  2253 => (x"f1",x"49",x"bf",x"d2"),
  2254 => (x"49",x"c0",x"87",x"fa"),
  2255 => (x"c2",x"87",x"da",x"f3"),
  2256 => (x"c0",x"48",x"f4",x"ce"),
  2257 => (x"f2",x"8e",x"f4",x"78"),
  2258 => (x"5e",x"0e",x"87",x"f4"),
  2259 => (x"0e",x"5d",x"5c",x"5b"),
  2260 => (x"c2",x"4c",x"71",x"1e"),
  2261 => (x"49",x"bf",x"ce",x"ee"),
  2262 => (x"4d",x"a1",x"cd",x"c1"),
  2263 => (x"69",x"81",x"d1",x"c1"),
  2264 => (x"02",x"9c",x"74",x"7e"),
  2265 => (x"a5",x"c4",x"87",x"cf"),
  2266 => (x"c2",x"7b",x"74",x"4b"),
  2267 => (x"49",x"bf",x"ce",x"ee"),
  2268 => (x"6e",x"87",x"d3",x"f2"),
  2269 => (x"05",x"9c",x"74",x"7b"),
  2270 => (x"4b",x"c0",x"87",x"c4"),
  2271 => (x"4b",x"c1",x"87",x"c2"),
  2272 => (x"d4",x"f2",x"49",x"73"),
  2273 => (x"02",x"66",x"d4",x"87"),
  2274 => (x"c0",x"49",x"87",x"c8"),
  2275 => (x"4a",x"70",x"87",x"ea"),
  2276 => (x"4a",x"c0",x"87",x"c2"),
  2277 => (x"5a",x"f8",x"ce",x"c2"),
  2278 => (x"87",x"e2",x"f1",x"26"),
  2279 => (x"14",x"11",x"12",x"58"),
  2280 => (x"23",x"1c",x"1b",x"1d"),
  2281 => (x"94",x"91",x"59",x"5a"),
  2282 => (x"f4",x"eb",x"f2",x"f5"),
  2283 => (x"00",x"00",x"00",x"00"),
  2284 => (x"00",x"00",x"00",x"00"),
  2285 => (x"00",x"00",x"00",x"00"),
  2286 => (x"ff",x"4a",x"71",x"1e"),
  2287 => (x"72",x"49",x"bf",x"c8"),
  2288 => (x"4f",x"26",x"48",x"a1"),
  2289 => (x"bf",x"c8",x"ff",x"1e"),
  2290 => (x"c0",x"c0",x"fe",x"89"),
  2291 => (x"a9",x"c0",x"c0",x"c0"),
  2292 => (x"c0",x"87",x"c4",x"01"),
  2293 => (x"c1",x"87",x"c2",x"4a"),
  2294 => (x"26",x"48",x"72",x"4a"),
  2295 => (x"5b",x"5e",x"0e",x"4f"),
  2296 => (x"71",x"0e",x"5d",x"5c"),
  2297 => (x"4c",x"d4",x"ff",x"4b"),
  2298 => (x"c0",x"48",x"66",x"d0"),
  2299 => (x"ff",x"49",x"d6",x"78"),
  2300 => (x"c3",x"87",x"e6",x"da"),
  2301 => (x"49",x"6c",x"7c",x"ff"),
  2302 => (x"71",x"99",x"ff",x"c3"),
  2303 => (x"f0",x"c3",x"49",x"4d"),
  2304 => (x"a9",x"e0",x"c1",x"99"),
  2305 => (x"c3",x"87",x"cb",x"05"),
  2306 => (x"48",x"6c",x"7c",x"ff"),
  2307 => (x"66",x"d0",x"98",x"c3"),
  2308 => (x"ff",x"c3",x"78",x"08"),
  2309 => (x"49",x"4a",x"6c",x"7c"),
  2310 => (x"ff",x"c3",x"31",x"c8"),
  2311 => (x"71",x"4a",x"6c",x"7c"),
  2312 => (x"c8",x"49",x"72",x"b2"),
  2313 => (x"7c",x"ff",x"c3",x"31"),
  2314 => (x"b2",x"71",x"4a",x"6c"),
  2315 => (x"31",x"c8",x"49",x"72"),
  2316 => (x"6c",x"7c",x"ff",x"c3"),
  2317 => (x"ff",x"b2",x"71",x"4a"),
  2318 => (x"e0",x"c0",x"48",x"d0"),
  2319 => (x"02",x"9b",x"73",x"78"),
  2320 => (x"7b",x"72",x"87",x"c2"),
  2321 => (x"4d",x"26",x"48",x"75"),
  2322 => (x"4b",x"26",x"4c",x"26"),
  2323 => (x"26",x"1e",x"4f",x"26"),
  2324 => (x"5b",x"5e",x"0e",x"4f"),
  2325 => (x"86",x"f8",x"0e",x"5c"),
  2326 => (x"a6",x"c8",x"1e",x"76"),
  2327 => (x"87",x"fd",x"fd",x"49"),
  2328 => (x"4b",x"70",x"86",x"c4"),
  2329 => (x"a8",x"c2",x"48",x"6e"),
  2330 => (x"87",x"f0",x"c2",x"03"),
  2331 => (x"f0",x"c3",x"4a",x"73"),
  2332 => (x"aa",x"d0",x"c1",x"9a"),
  2333 => (x"c1",x"87",x"c7",x"02"),
  2334 => (x"c2",x"05",x"aa",x"e0"),
  2335 => (x"49",x"73",x"87",x"de"),
  2336 => (x"c3",x"02",x"99",x"c8"),
  2337 => (x"87",x"c6",x"ff",x"87"),
  2338 => (x"9c",x"c3",x"4c",x"73"),
  2339 => (x"c1",x"05",x"ac",x"c2"),
  2340 => (x"66",x"c4",x"87",x"c2"),
  2341 => (x"71",x"31",x"c9",x"49"),
  2342 => (x"4a",x"66",x"c4",x"1e"),
  2343 => (x"ee",x"c2",x"92",x"d4"),
  2344 => (x"81",x"72",x"49",x"d6"),
  2345 => (x"87",x"c7",x"d4",x"fe"),
  2346 => (x"d7",x"ff",x"49",x"d8"),
  2347 => (x"c0",x"c8",x"87",x"eb"),
  2348 => (x"c6",x"dd",x"c2",x"1e"),
  2349 => (x"e2",x"f0",x"fd",x"49"),
  2350 => (x"48",x"d0",x"ff",x"87"),
  2351 => (x"c2",x"78",x"e0",x"c0"),
  2352 => (x"cc",x"1e",x"c6",x"dd"),
  2353 => (x"92",x"d4",x"4a",x"66"),
  2354 => (x"49",x"d6",x"ee",x"c2"),
  2355 => (x"d2",x"fe",x"81",x"72"),
  2356 => (x"86",x"cc",x"87",x"da"),
  2357 => (x"c1",x"05",x"ac",x"c1"),
  2358 => (x"66",x"c4",x"87",x"c2"),
  2359 => (x"71",x"31",x"c9",x"49"),
  2360 => (x"4a",x"66",x"c4",x"1e"),
  2361 => (x"ee",x"c2",x"92",x"d4"),
  2362 => (x"81",x"72",x"49",x"d6"),
  2363 => (x"87",x"ff",x"d2",x"fe"),
  2364 => (x"1e",x"c6",x"dd",x"c2"),
  2365 => (x"d4",x"4a",x"66",x"c8"),
  2366 => (x"d6",x"ee",x"c2",x"92"),
  2367 => (x"fe",x"81",x"72",x"49"),
  2368 => (x"d7",x"87",x"e6",x"d0"),
  2369 => (x"d0",x"d6",x"ff",x"49"),
  2370 => (x"1e",x"c0",x"c8",x"87"),
  2371 => (x"49",x"c6",x"dd",x"c2"),
  2372 => (x"87",x"f1",x"ee",x"fd"),
  2373 => (x"d0",x"ff",x"86",x"cc"),
  2374 => (x"78",x"e0",x"c0",x"48"),
  2375 => (x"e7",x"fc",x"8e",x"f8"),
  2376 => (x"5b",x"5e",x"0e",x"87"),
  2377 => (x"1e",x"0e",x"5d",x"5c"),
  2378 => (x"d4",x"ff",x"4d",x"71"),
  2379 => (x"7e",x"66",x"d4",x"4c"),
  2380 => (x"a8",x"b7",x"c3",x"48"),
  2381 => (x"c0",x"87",x"c5",x"06"),
  2382 => (x"87",x"e2",x"c1",x"48"),
  2383 => (x"e0",x"fe",x"49",x"75"),
  2384 => (x"1e",x"75",x"87",x"fe"),
  2385 => (x"d4",x"4b",x"66",x"c4"),
  2386 => (x"d6",x"ee",x"c2",x"93"),
  2387 => (x"fe",x"49",x"73",x"83"),
  2388 => (x"c8",x"87",x"fa",x"cb"),
  2389 => (x"ff",x"4b",x"6b",x"83"),
  2390 => (x"e1",x"c8",x"48",x"d0"),
  2391 => (x"73",x"7c",x"dd",x"78"),
  2392 => (x"99",x"ff",x"c3",x"49"),
  2393 => (x"49",x"73",x"7c",x"71"),
  2394 => (x"c3",x"29",x"b7",x"c8"),
  2395 => (x"7c",x"71",x"99",x"ff"),
  2396 => (x"b7",x"d0",x"49",x"73"),
  2397 => (x"99",x"ff",x"c3",x"29"),
  2398 => (x"49",x"73",x"7c",x"71"),
  2399 => (x"71",x"29",x"b7",x"d8"),
  2400 => (x"7c",x"7c",x"c0",x"7c"),
  2401 => (x"7c",x"7c",x"7c",x"7c"),
  2402 => (x"7c",x"7c",x"7c",x"7c"),
  2403 => (x"e0",x"c0",x"7c",x"7c"),
  2404 => (x"1e",x"66",x"c4",x"78"),
  2405 => (x"d4",x"ff",x"49",x"dc"),
  2406 => (x"86",x"c8",x"87",x"e4"),
  2407 => (x"fa",x"26",x"48",x"73"),
  2408 => (x"5e",x"0e",x"87",x"e4"),
  2409 => (x"0e",x"5d",x"5c",x"5b"),
  2410 => (x"ff",x"7e",x"71",x"1e"),
  2411 => (x"1e",x"6e",x"4b",x"d4"),
  2412 => (x"49",x"fe",x"ee",x"c2"),
  2413 => (x"87",x"d5",x"ca",x"fe"),
  2414 => (x"4d",x"70",x"86",x"c4"),
  2415 => (x"c3",x"c3",x"02",x"9d"),
  2416 => (x"c6",x"ef",x"c2",x"87"),
  2417 => (x"49",x"6e",x"4c",x"bf"),
  2418 => (x"87",x"f4",x"de",x"fe"),
  2419 => (x"c8",x"48",x"d0",x"ff"),
  2420 => (x"d6",x"c1",x"78",x"c5"),
  2421 => (x"15",x"4a",x"c0",x"7b"),
  2422 => (x"c0",x"82",x"c1",x"7b"),
  2423 => (x"04",x"aa",x"b7",x"e0"),
  2424 => (x"d0",x"ff",x"87",x"f5"),
  2425 => (x"c8",x"78",x"c4",x"48"),
  2426 => (x"d3",x"c1",x"78",x"c5"),
  2427 => (x"c4",x"7b",x"c1",x"7b"),
  2428 => (x"02",x"9c",x"74",x"78"),
  2429 => (x"c2",x"87",x"fc",x"c1"),
  2430 => (x"c8",x"7e",x"c6",x"dd"),
  2431 => (x"c0",x"8c",x"4d",x"c0"),
  2432 => (x"c6",x"03",x"ac",x"b7"),
  2433 => (x"a4",x"c0",x"c8",x"87"),
  2434 => (x"c2",x"4c",x"c0",x"4d"),
  2435 => (x"bf",x"97",x"f7",x"e9"),
  2436 => (x"02",x"99",x"d0",x"49"),
  2437 => (x"1e",x"c0",x"87",x"d2"),
  2438 => (x"49",x"fe",x"ee",x"c2"),
  2439 => (x"87",x"c9",x"cc",x"fe"),
  2440 => (x"49",x"70",x"86",x"c4"),
  2441 => (x"87",x"ef",x"c0",x"4a"),
  2442 => (x"1e",x"c6",x"dd",x"c2"),
  2443 => (x"49",x"fe",x"ee",x"c2"),
  2444 => (x"87",x"f5",x"cb",x"fe"),
  2445 => (x"49",x"70",x"86",x"c4"),
  2446 => (x"48",x"d0",x"ff",x"4a"),
  2447 => (x"c1",x"78",x"c5",x"c8"),
  2448 => (x"97",x"6e",x"7b",x"d4"),
  2449 => (x"48",x"6e",x"7b",x"bf"),
  2450 => (x"7e",x"70",x"80",x"c1"),
  2451 => (x"ff",x"05",x"8d",x"c1"),
  2452 => (x"d0",x"ff",x"87",x"f0"),
  2453 => (x"72",x"78",x"c4",x"48"),
  2454 => (x"87",x"c5",x"05",x"9a"),
  2455 => (x"e5",x"c0",x"48",x"c0"),
  2456 => (x"c2",x"1e",x"c1",x"87"),
  2457 => (x"fe",x"49",x"fe",x"ee"),
  2458 => (x"c4",x"87",x"dd",x"c9"),
  2459 => (x"05",x"9c",x"74",x"86"),
  2460 => (x"ff",x"87",x"c4",x"fe"),
  2461 => (x"c5",x"c8",x"48",x"d0"),
  2462 => (x"7b",x"d3",x"c1",x"78"),
  2463 => (x"78",x"c4",x"7b",x"c0"),
  2464 => (x"87",x"c2",x"48",x"c1"),
  2465 => (x"26",x"26",x"48",x"c0"),
  2466 => (x"26",x"4c",x"26",x"4d"),
  2467 => (x"0e",x"4f",x"26",x"4b"),
  2468 => (x"0e",x"5c",x"5b",x"5e"),
  2469 => (x"66",x"cc",x"4b",x"71"),
  2470 => (x"4c",x"87",x"d8",x"02"),
  2471 => (x"02",x"8c",x"f0",x"c0"),
  2472 => (x"4a",x"74",x"87",x"d8"),
  2473 => (x"d1",x"02",x"8a",x"c1"),
  2474 => (x"cd",x"02",x"8a",x"87"),
  2475 => (x"c9",x"02",x"8a",x"87"),
  2476 => (x"73",x"87",x"d7",x"87"),
  2477 => (x"87",x"ea",x"fb",x"49"),
  2478 => (x"1e",x"74",x"87",x"d0"),
  2479 => (x"e0",x"f9",x"49",x"c0"),
  2480 => (x"73",x"1e",x"74",x"87"),
  2481 => (x"87",x"d9",x"f9",x"49"),
  2482 => (x"fc",x"fe",x"86",x"c8"),
  2483 => (x"c2",x"1e",x"00",x"87"),
  2484 => (x"49",x"bf",x"dc",x"dc"),
  2485 => (x"dc",x"c2",x"b9",x"c1"),
  2486 => (x"d4",x"ff",x"59",x"e0"),
  2487 => (x"78",x"ff",x"c3",x"48"),
  2488 => (x"c8",x"48",x"d0",x"ff"),
  2489 => (x"d4",x"ff",x"78",x"e1"),
  2490 => (x"c4",x"78",x"c1",x"48"),
  2491 => (x"ff",x"78",x"71",x"31"),
  2492 => (x"e0",x"c0",x"48",x"d0"),
  2493 => (x"1e",x"4f",x"26",x"78"),
  2494 => (x"1e",x"d0",x"dc",x"c2"),
  2495 => (x"49",x"fe",x"ee",x"c2"),
  2496 => (x"87",x"c9",x"c5",x"fe"),
  2497 => (x"98",x"70",x"86",x"c4"),
  2498 => (x"ff",x"87",x"c3",x"02"),
  2499 => (x"4f",x"26",x"87",x"c0"),
  2500 => (x"48",x"4b",x"35",x"31"),
  2501 => (x"20",x"20",x"20",x"5a"),
  2502 => (x"00",x"47",x"46",x"43"),
  2503 => (x"00",x"00",x"00",x"00"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

