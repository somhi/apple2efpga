library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom2 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"01010000",
     1 => x"01017f7f",
     2 => x"7f3f0000",
     3 => x"3f7f4040",
     4 => x"3f0f0000",
     5 => x"0f3f7070",
     6 => x"307f7f00",
     7 => x"7f7f3018",
     8 => x"36634100",
     9 => x"63361c1c",
    10 => x"06030141",
    11 => x"03067c7c",
    12 => x"59716101",
    13 => x"4143474d",
    14 => x"7f000000",
    15 => x"0041417f",
    16 => x"06030100",
    17 => x"6030180c",
    18 => x"41000040",
    19 => x"007f7f41",
    20 => x"060c0800",
    21 => x"080c0603",
    22 => x"80808000",
    23 => x"80808080",
    24 => x"00000000",
    25 => x"00040703",
    26 => x"74200000",
    27 => x"787c5454",
    28 => x"7f7f0000",
    29 => x"387c4444",
    30 => x"7c380000",
    31 => x"00444444",
    32 => x"7c380000",
    33 => x"7f7f4444",
    34 => x"7c380000",
    35 => x"185c5454",
    36 => x"7e040000",
    37 => x"0005057f",
    38 => x"bc180000",
    39 => x"7cfca4a4",
    40 => x"7f7f0000",
    41 => x"787c0404",
    42 => x"00000000",
    43 => x"00407d3d",
    44 => x"80800000",
    45 => x"007dfd80",
    46 => x"7f7f0000",
    47 => x"446c3810",
    48 => x"00000000",
    49 => x"00407f3f",
    50 => x"0c7c7c00",
    51 => x"787c0c18",
    52 => x"7c7c0000",
    53 => x"787c0404",
    54 => x"7c380000",
    55 => x"387c4444",
    56 => x"fcfc0000",
    57 => x"183c2424",
    58 => x"3c180000",
    59 => x"fcfc2424",
    60 => x"7c7c0000",
    61 => x"080c0404",
    62 => x"5c480000",
    63 => x"20745454",
    64 => x"3f040000",
    65 => x"0044447f",
    66 => x"7c3c0000",
    67 => x"7c7c4040",
    68 => x"3c1c0000",
    69 => x"1c3c6060",
    70 => x"607c3c00",
    71 => x"3c7c6030",
    72 => x"386c4400",
    73 => x"446c3810",
    74 => x"bc1c0000",
    75 => x"1c3c60e0",
    76 => x"64440000",
    77 => x"444c5c74",
    78 => x"08080000",
    79 => x"4141773e",
    80 => x"00000000",
    81 => x"00007f7f",
    82 => x"41410000",
    83 => x"08083e77",
    84 => x"01010200",
    85 => x"01020203",
    86 => x"7f7f7f00",
    87 => x"7f7f7f7f",
    88 => x"1c080800",
    89 => x"7f3e3e1c",
    90 => x"3e7f7f7f",
    91 => x"081c1c3e",
    92 => x"18100008",
    93 => x"10187c7c",
    94 => x"30100000",
    95 => x"10307c7c",
    96 => x"60301000",
    97 => x"061e7860",
    98 => x"3c664200",
    99 => x"42663c18",
   100 => x"6a387800",
   101 => x"386cc6c2",
   102 => x"00006000",
   103 => x"60000060",
   104 => x"5b5e0e00",
   105 => x"1e0e5d5c",
   106 => x"cbc34c71",
   107 => x"c04dbfce",
   108 => x"741ec04b",
   109 => x"87c702ab",
   110 => x"c048a6c4",
   111 => x"c487c578",
   112 => x"78c148a6",
   113 => x"731e66c4",
   114 => x"87dfee49",
   115 => x"e0c086c8",
   116 => x"87efef49",
   117 => x"6a4aa5c4",
   118 => x"87f0f049",
   119 => x"cb87c6f1",
   120 => x"c883c185",
   121 => x"ff04abb7",
   122 => x"262687c7",
   123 => x"264c264d",
   124 => x"1e4f264b",
   125 => x"cbc34a71",
   126 => x"cbc35ad2",
   127 => x"78c748d2",
   128 => x"87ddfe49",
   129 => x"731e4f26",
   130 => x"c04a711e",
   131 => x"d303aab7",
   132 => x"cdd5c287",
   133 => x"87c405bf",
   134 => x"87c24bc1",
   135 => x"d5c24bc0",
   136 => x"87c45bd1",
   137 => x"5ad1d5c2",
   138 => x"bfcdd5c2",
   139 => x"c19ac14a",
   140 => x"ec49a2c0",
   141 => x"48fc87e8",
   142 => x"bfcdd5c2",
   143 => x"87effe78",
   144 => x"cdd5c21e",
   145 => x"e7c049bf",
   146 => x"cbc387e4",
   147 => x"bfe848c6",
   148 => x"c2cbc378",
   149 => x"78bfec48",
   150 => x"bfc6cbc3",
   151 => x"ffc3494a",
   152 => x"2ab7c899",
   153 => x"b0714872",
   154 => x"58cecbc3",
   155 => x"5e0e4f26",
   156 => x"0e5d5c5b",
   157 => x"c7ff4b71",
   158 => x"c1cbc387",
   159 => x"7350c048",
   160 => x"87d3e549",
   161 => x"c24c4970",
   162 => x"49eecb9c",
   163 => x"7087c6cb",
   164 => x"cbc34d49",
   165 => x"05bf97c1",
   166 => x"d087e2c1",
   167 => x"cbc34966",
   168 => x"0599bfca",
   169 => x"66d487d6",
   170 => x"c2cbc349",
   171 => x"cb0599bf",
   172 => x"e4497387",
   173 => x"987087e1",
   174 => x"87c1c102",
   175 => x"fffd4cc1",
   176 => x"ca497587",
   177 => x"987087db",
   178 => x"c387c602",
   179 => x"c148c1cb",
   180 => x"c1cbc350",
   181 => x"c005bf97",
   182 => x"cbc387e3",
   183 => x"d049bfca",
   184 => x"ff059966",
   185 => x"cbc387d6",
   186 => x"d449bfc2",
   187 => x"ff059966",
   188 => x"497387ca",
   189 => x"7087e0e3",
   190 => x"fffe0598",
   191 => x"fb487487",
   192 => x"5e0e87e9",
   193 => x"0e5d5c5b",
   194 => x"4dc086f4",
   195 => x"7ebfec4c",
   196 => x"c348a6c4",
   197 => x"78bfcecb",
   198 => x"1ec01ec1",
   199 => x"cdfd49c7",
   200 => x"7086c887",
   201 => x"87cd0298",
   202 => x"d9fb49ff",
   203 => x"49dac187",
   204 => x"c187e4e2",
   205 => x"c1cbc34d",
   206 => x"c302bf97",
   207 => x"87c6d587",
   208 => x"bfc6cbc3",
   209 => x"cdd5c24b",
   210 => x"ebc005bf",
   211 => x"49fdc387",
   212 => x"c387c4e2",
   213 => x"fee149fa",
   214 => x"c3497387",
   215 => x"1e7199ff",
   216 => x"e4c049c0",
   217 => x"497387ec",
   218 => x"7129b7c8",
   219 => x"c049c11e",
   220 => x"c887dfe4",
   221 => x"87fbc586",
   222 => x"bfcacbc3",
   223 => x"dd029b4b",
   224 => x"c9d5c287",
   225 => x"d8c749bf",
   226 => x"05987087",
   227 => x"4bc087c4",
   228 => x"e0c287d2",
   229 => x"87fdc649",
   230 => x"58cdd5c2",
   231 => x"d5c287c6",
   232 => x"78c048c9",
   233 => x"99c24973",
   234 => x"c387cd05",
   235 => x"e6e049eb",
   236 => x"c2497087",
   237 => x"87c20299",
   238 => x"49734cfb",
   239 => x"cd0599c1",
   240 => x"49f4c387",
   241 => x"7087d0e0",
   242 => x"0299c249",
   243 => x"4cfa87c2",
   244 => x"99c84973",
   245 => x"c387ce05",
   246 => x"dfff49f5",
   247 => x"497087f9",
   248 => x"d40299c2",
   249 => x"d2cbc387",
   250 => x"87c902bf",
   251 => x"c388c148",
   252 => x"c258d6cb",
   253 => x"c14cff87",
   254 => x"c449734d",
   255 => x"87ce0599",
   256 => x"ff49f2c3",
   257 => x"7087d0df",
   258 => x"0299c249",
   259 => x"cbc387db",
   260 => x"487ebfd2",
   261 => x"03a8b7c7",
   262 => x"486e87cb",
   263 => x"cbc380c1",
   264 => x"c2c058d6",
   265 => x"c14cfe87",
   266 => x"49fdc34d",
   267 => x"87e7deff",
   268 => x"99c24970",
   269 => x"c387d502",
   270 => x"02bfd2cb",
   271 => x"c387c9c0",
   272 => x"c048d2cb",
   273 => x"87c2c078",
   274 => x"4dc14cfd",
   275 => x"ff49fac3",
   276 => x"7087c4de",
   277 => x"0299c249",
   278 => x"cbc387d9",
   279 => x"c748bfd2",
   280 => x"c003a8b7",
   281 => x"cbc387c9",
   282 => x"78c748d2",
   283 => x"fc87c2c0",
   284 => x"c04dc14c",
   285 => x"c003acb7",
   286 => x"66c487d1",
   287 => x"82d8c14a",
   288 => x"c6c0026a",
   289 => x"744b6a87",
   290 => x"c00f7349",
   291 => x"1ef0c31e",
   292 => x"f749dac1",
   293 => x"86c887d8",
   294 => x"c0029870",
   295 => x"a6c887e2",
   296 => x"d2cbc348",
   297 => x"66c878bf",
   298 => x"c491cb49",
   299 => x"80714866",
   300 => x"bf6e7e70",
   301 => x"87c8c002",
   302 => x"c84bbf6e",
   303 => x"0f734966",
   304 => x"c0029d75",
   305 => x"cbc387c8",
   306 => x"f349bfd2",
   307 => x"d5c287d3",
   308 => x"c002bfd1",
   309 => x"c24987dd",
   310 => x"987087c7",
   311 => x"87d3c002",
   312 => x"bfd2cbc3",
   313 => x"87f9f249",
   314 => x"d9f449c0",
   315 => x"d1d5c287",
   316 => x"f478c048",
   317 => x"87f3f38e",
   318 => x"5c5b5e0e",
   319 => x"711e0e5d",
   320 => x"cecbc34c",
   321 => x"cdc149bf",
   322 => x"d1c14da1",
   323 => x"747e6981",
   324 => x"87cf029c",
   325 => x"744ba5c4",
   326 => x"cecbc37b",
   327 => x"d2f349bf",
   328 => x"747b6e87",
   329 => x"87c4059c",
   330 => x"87c24bc0",
   331 => x"49734bc1",
   332 => x"d487d3f3",
   333 => x"87c70266",
   334 => x"7087da49",
   335 => x"c087c24a",
   336 => x"d5d5c24a",
   337 => x"e2f2265a",
   338 => x"00000087",
   339 => x"00000000",
   340 => x"00000000",
   341 => x"4a711e00",
   342 => x"49bfc8ff",
   343 => x"2648a172",
   344 => x"c8ff1e4f",
   345 => x"c0fe89bf",
   346 => x"c0c0c0c0",
   347 => x"87c401a9",
   348 => x"87c24ac0",
   349 => x"48724ac1",
   350 => x"5e0e4f26",
   351 => x"0e5d5c5b",
   352 => x"d4ff4b71",
   353 => x"4866d04c",
   354 => x"49d678c0",
   355 => x"87c7dbff",
   356 => x"6c7cffc3",
   357 => x"99ffc349",
   358 => x"c3494d71",
   359 => x"e0c199f0",
   360 => x"87cb05a9",
   361 => x"6c7cffc3",
   362 => x"d098c348",
   363 => x"c3780866",
   364 => x"4a6c7cff",
   365 => x"c331c849",
   366 => x"4a6c7cff",
   367 => x"4972b271",
   368 => x"ffc331c8",
   369 => x"714a6c7c",
   370 => x"c84972b2",
   371 => x"7cffc331",
   372 => x"b2714a6c",
   373 => x"c048d0ff",
   374 => x"9b7378e0",
   375 => x"7287c202",
   376 => x"2648757b",
   377 => x"264c264d",
   378 => x"1e4f264b",
   379 => x"5e0e4f26",
   380 => x"f80e5c5b",
   381 => x"c81e7686",
   382 => x"fdfd49a6",
   383 => x"7086c487",
   384 => x"c2486e4b",
   385 => x"cac303a8",
   386 => x"c34a7387",
   387 => x"d0c19af0",
   388 => x"87c702aa",
   389 => x"05aae0c1",
   390 => x"7387f8c2",
   391 => x"0299c849",
   392 => x"c6ff87c3",
   393 => x"c34c7387",
   394 => x"05acc29c",
   395 => x"c487cfc1",
   396 => x"31c94966",
   397 => x"66c41e71",
   398 => x"92d8c24a",
   399 => x"49d6cbc3",
   400 => x"d3fe8172",
   401 => x"66c487c0",
   402 => x"e3c01e49",
   403 => x"ebd8ff49",
   404 => x"ff49d887",
   405 => x"c887c0d8",
   406 => x"fac21ec0",
   407 => x"ebfd49c6",
   408 => x"d0ff87de",
   409 => x"78e0c048",
   410 => x"1ec6fac2",
   411 => x"c24a66d0",
   412 => x"cbc392d8",
   413 => x"817249d6",
   414 => x"87c8cefe",
   415 => x"acc186d0",
   416 => x"87cfc105",
   417 => x"c94966c4",
   418 => x"c41e7131",
   419 => x"d8c24a66",
   420 => x"d6cbc392",
   421 => x"fe817249",
   422 => x"c287ebd1",
   423 => x"c81ec6fa",
   424 => x"d8c24a66",
   425 => x"d6cbc392",
   426 => x"fe817249",
   427 => x"c887d2cc",
   428 => x"c01e4966",
   429 => x"d7ff49e3",
   430 => x"49d787c2",
   431 => x"87d7d6ff",
   432 => x"c21ec0c8",
   433 => x"fd49c6fa",
   434 => x"d087dfe9",
   435 => x"48d0ff86",
   436 => x"f878e0c0",
   437 => x"87cdfc8e",
   438 => x"5c5b5e0e",
   439 => x"711e0e5d",
   440 => x"4cd4ff4d",
   441 => x"487e66d4",
   442 => x"06a8b7c3",
   443 => x"48c087c5",
   444 => x"7587e3c1",
   445 => x"f4e1fe49",
   446 => x"c41e7587",
   447 => x"d8c24b66",
   448 => x"d6cbc393",
   449 => x"fe497383",
   450 => x"c887e9c6",
   451 => x"ff4b6b83",
   452 => x"e1c848d0",
   453 => x"737cdd78",
   454 => x"99ffc349",
   455 => x"49737c71",
   456 => x"c329b7c8",
   457 => x"7c7199ff",
   458 => x"b7d04973",
   459 => x"99ffc329",
   460 => x"49737c71",
   461 => x"7129b7d8",
   462 => x"7c7cc07c",
   463 => x"7c7c7c7c",
   464 => x"7c7c7c7c",
   465 => x"e0c07c7c",
   466 => x"1e66c478",
   467 => x"d4ff49dc",
   468 => x"86c887ea",
   469 => x"fa264873",
   470 => x"5e0e87c9",
   471 => x"0e5d5c5b",
   472 => x"ff7e711e",
   473 => x"1e6e4bd4",
   474 => x"49c6d0c3",
   475 => x"87c4c5fe",
   476 => x"4d7086c4",
   477 => x"c3c3029d",
   478 => x"ced0c387",
   479 => x"496e4cbf",
   480 => x"87e9dffe",
   481 => x"c848d0ff",
   482 => x"d6c178c5",
   483 => x"154ac07b",
   484 => x"c082c17b",
   485 => x"04aab7e0",
   486 => x"d0ff87f5",
   487 => x"c878c448",
   488 => x"d3c178c5",
   489 => x"c47bc17b",
   490 => x"029c7478",
   491 => x"c287fcc1",
   492 => x"c87ec6fa",
   493 => x"c08c4dc0",
   494 => x"c603acb7",
   495 => x"a4c0c887",
   496 => x"c34cc04d",
   497 => x"bf97f7c6",
   498 => x"0299d049",
   499 => x"1ec087d2",
   500 => x"49c6d0c3",
   501 => x"87e9c7fe",
   502 => x"497086c4",
   503 => x"87efc04a",
   504 => x"1ec6fac2",
   505 => x"49c6d0c3",
   506 => x"87d5c7fe",
   507 => x"497086c4",
   508 => x"48d0ff4a",
   509 => x"c178c5c8",
   510 => x"976e7bd4",
   511 => x"486e7bbf",
   512 => x"7e7080c1",
   513 => x"ff058dc1",
   514 => x"d0ff87f0",
   515 => x"7278c448",
   516 => x"87c5059a",
   517 => x"e5c048c0",
   518 => x"c31ec187",
   519 => x"fe49c6d0",
   520 => x"c487fdc4",
   521 => x"059c7486",
   522 => x"ff87c4fe",
   523 => x"c5c848d0",
   524 => x"7bd3c178",
   525 => x"78c47bc0",
   526 => x"87c248c1",
   527 => x"262648c0",
   528 => x"264c264d",
   529 => x"0e4f264b",
   530 => x"0e5c5b5e",
   531 => x"66cc4b71",
   532 => x"4c87d802",
   533 => x"028cf0c0",
   534 => x"4a7487d8",
   535 => x"d1028ac1",
   536 => x"cd028a87",
   537 => x"c9028a87",
   538 => x"7387d787",
   539 => x"87eafb49",
   540 => x"1e7487d0",
   541 => x"dff949c0",
   542 => x"731e7487",
   543 => x"87d8f949",
   544 => x"fcfe86c8",
   545 => x"c21e0087",
   546 => x"49bfefe2",
   547 => x"e2c2b9c1",
   548 => x"d4ff59f3",
   549 => x"78ffc348",
   550 => x"c848d0ff",
   551 => x"d4ff78e1",
   552 => x"c478c148",
   553 => x"ff787131",
   554 => x"e0c048d0",
   555 => x"004f2678",
   556 => x"1e000000",
   557 => x"87edc3ff",
   558 => x"c24966c4",
   559 => x"cd0299c0",
   560 => x"1ee0c387",
   561 => x"49e3cac3",
   562 => x"87fcc4ff",
   563 => x"66c486c4",
   564 => x"99c0c449",
   565 => x"c387cd02",
   566 => x"cac31ef0",
   567 => x"c4ff49e3",
   568 => x"86c487e6",
   569 => x"c14966c4",
   570 => x"1e7199ff",
   571 => x"49e3cac3",
   572 => x"87d4c4ff",
   573 => x"87e5c2ff",
   574 => x"0e4f2626",
   575 => x"5d5c5b5e",
   576 => x"86dcff0e",
   577 => x"d2c37ec0",
   578 => x"c249bfe2",
   579 => x"721e7181",
   580 => x"fd4ac61e",
   581 => x"7187e2df",
   582 => x"264a2648",
   583 => x"58a6c849",
   584 => x"bfe2d2c3",
   585 => x"7181c449",
   586 => x"c61e721e",
   587 => x"c8dffd4a",
   588 => x"26487187",
   589 => x"cc49264a",
   590 => x"4cc058a6",
   591 => x"91c44974",
   592 => x"6981d0fe",
   593 => x"c349744a",
   594 => x"81bfe2d2",
   595 => x"d2c391c4",
   596 => x"797281f2",
   597 => x"87d1029a",
   598 => x"89c14972",
   599 => x"486e9a71",
   600 => x"7e7080c1",
   601 => x"ef059a72",
   602 => x"c284c187",
   603 => x"ff04acb7",
   604 => x"486e87ca",
   605 => x"a8b7fcc0",
   606 => x"87ffc804",
   607 => x"4a744cc0",
   608 => x"c48266c4",
   609 => x"f2d2c392",
   610 => x"c8497482",
   611 => x"91c48166",
   612 => x"81f2d2c3",
   613 => x"49694a6a",
   614 => x"4b74b972",
   615 => x"bfe2d2c3",
   616 => x"c393c483",
   617 => x"6b83f2d2",
   618 => x"714872ba",
   619 => x"58a6d098",
   620 => x"d2c34974",
   621 => x"c481bfe2",
   622 => x"f2d2c391",
   623 => x"d07e6981",
   624 => x"78c048a6",
   625 => x"df4966cc",
   626 => x"c0c70229",
   627 => x"c04a7487",
   628 => x"66d092e0",
   629 => x"48ffc082",
   630 => x"4a708872",
   631 => x"c048a6d4",
   632 => x"c080c478",
   633 => x"df496e78",
   634 => x"a6e0c029",
   635 => x"ded2c359",
   636 => x"7278c148",
   637 => x"b731c349",
   638 => x"c0b1722a",
   639 => x"91c499ff",
   640 => x"4dd9f5c2",
   641 => x"4b6d8571",
   642 => x"c0c0c449",
   643 => x"f3c00299",
   644 => x"0266dc87",
   645 => x"80c887c8",
   646 => x"c57840c0",
   647 => x"d2c387ef",
   648 => x"78c148e6",
   649 => x"bfead2c3",
   650 => x"87e1c505",
   651 => x"f81ed8c1",
   652 => x"fef949a0",
   653 => x"1ed8c587",
   654 => x"49ded2c3",
   655 => x"c887f4f9",
   656 => x"87c9c586",
   657 => x"d80266dc",
   658 => x"c2497387",
   659 => x"0299c0c0",
   660 => x"d087c3c0",
   661 => x"486d2bb7",
   662 => x"98fffffd",
   663 => x"fac07d70",
   664 => x"e6d2c387",
   665 => x"f2c002bf",
   666 => x"d0487387",
   667 => x"e4c028b7",
   668 => x"987058a6",
   669 => x"87e3c002",
   670 => x"bfeed2c3",
   671 => x"c0e0c049",
   672 => x"cac00299",
   673 => x"c0497087",
   674 => x"0299c0e0",
   675 => x"6d87ccc0",
   676 => x"c0c0c248",
   677 => x"c07d70b0",
   678 => x"734b66e0",
   679 => x"c0c0c849",
   680 => x"c7c20299",
   681 => x"eed2c387",
   682 => x"c0cc4abf",
   683 => x"cfc0029a",
   684 => x"8ac0c487",
   685 => x"87d8c002",
   686 => x"f9c0028a",
   687 => x"87ddc187",
   688 => x"ffc34973",
   689 => x"c291c299",
   690 => x"1181cdf5",
   691 => x"87dcc14b",
   692 => x"ffc34973",
   693 => x"c291c299",
   694 => x"c181cdf5",
   695 => x"dc4b1181",
   696 => x"c8c00266",
   697 => x"48a6d887",
   698 => x"ffc078d2",
   699 => x"48a6d487",
   700 => x"c078d2c4",
   701 => x"497387f6",
   702 => x"c299ffc3",
   703 => x"cdf5c291",
   704 => x"1181c181",
   705 => x"0266dc4b",
   706 => x"d887c9c0",
   707 => x"d9c148a6",
   708 => x"87d8c078",
   709 => x"c548a6d4",
   710 => x"cfc078d9",
   711 => x"c3497387",
   712 => x"91c299ff",
   713 => x"81cdf5c2",
   714 => x"4b1181c1",
   715 => x"c00266dc",
   716 => x"497387dc",
   717 => x"fcc7b9ff",
   718 => x"487199c0",
   719 => x"bfeed2c3",
   720 => x"f2d2c398",
   721 => x"9bffc358",
   722 => x"c0b3c0c4",
   723 => x"497387d4",
   724 => x"99c0fcc7",
   725 => x"d2c34871",
   726 => x"c3b0bfee",
   727 => x"c358f2d2",
   728 => x"66d49bff",
   729 => x"87cac002",
   730 => x"ded2c31e",
   731 => x"87c3f549",
   732 => x"1e7386c4",
   733 => x"49ded2c3",
   734 => x"c487f8f4",
   735 => x"0266d886",
   736 => x"1e87cac0",
   737 => x"49ded2c3",
   738 => x"c487e8f4",
   739 => x"4866cc86",
   740 => x"a6d030c1",
   741 => x"c1486e58",
   742 => x"d07e7030",
   743 => x"80c14866",
   744 => x"c058a6d4",
   745 => x"04a8b7e0",
   746 => x"c187d9f8",
   747 => x"acb7c284",
   748 => x"87caf704",
   749 => x"48e2d2c3",
   750 => x"ff7866c4",
   751 => x"4d268edc",
   752 => x"4b264c26",
   753 => x"c01e4f26",
   754 => x"c449724a",
   755 => x"f2d2c391",
   756 => x"c179ff81",
   757 => x"aab7c682",
   758 => x"c387ee04",
   759 => x"c048e2d2",
   760 => x"80c87840",
   761 => x"4f2678c0",
   762 => x"711e731e",
   763 => x"c1cbc34b",
   764 => x"c002bf97",
   765 => x"497387e9",
   766 => x"e4c191cb",
   767 => x"81ca81dc",
   768 => x"99496997",
   769 => x"c287d805",
   770 => x"c71ec11e",
   771 => x"fec3ff49",
   772 => x"c11ec287",
   773 => x"ff49c71e",
   774 => x"d087f4c3",
   775 => x"7387cc86",
   776 => x"c1dcfe49",
   777 => x"fe497387",
   778 => x"fe87fbdb",
   779 => x"731e87d4",
   780 => x"f34b711e",
   781 => x"497387c5",
   782 => x"87fdfafe",
   783 => x"0e87c3fe",
   784 => x"5d5c5b5e",
   785 => x"6b4b710e",
   786 => x"c0c4f84a",
   787 => x"c0fcc74d",
   788 => x"4966d04c",
   789 => x"cf0299c2",
   790 => x"4966d487",
   791 => x"718909c0",
   792 => x"d434c44c",
   793 => x"87d78a66",
   794 => x"c14966d0",
   795 => x"87ca0299",
   796 => x"c44d66d4",
   797 => x"8266d435",
   798 => x"92cf87c5",
   799 => x"752ab7c4",
   800 => x"c103aab7",
   801 => x"b7744a87",
   802 => x"87c106aa",
   803 => x"fc7b724a",
   804 => x"5e0e87ec",
   805 => x"710e5c5b",
   806 => x"4abfec4c",
   807 => x"fcfe49c5",
   808 => x"987087f5",
   809 => x"c287c702",
   810 => x"df48d9f9",
   811 => x"49c678f0",
   812 => x"87e3fcfe",
   813 => x"c7029870",
   814 => x"d9f9c287",
   815 => x"78c0cc48",
   816 => x"fcfe49c4",
   817 => x"987087d1",
   818 => x"c287c702",
   819 => x"c448d9f9",
   820 => x"49cc78c0",
   821 => x"87fffbfe",
   822 => x"c7029870",
   823 => x"d9f9c287",
   824 => x"78c0c148",
   825 => x"741e66cc",
   826 => x"e4fefe49",
   827 => x"d9f9c287",
   828 => x"66d41ebf",
   829 => x"c24b741e",
   830 => x"c84a7493",
   831 => x"e2d3c392",
   832 => x"fc817249",
   833 => x"f9c287f9",
   834 => x"dc1ebfd9",
   835 => x"b7c24966",
   836 => x"731e7129",
   837 => x"c392c44a",
   838 => x"7249e6d3",
   839 => x"87dffc81",
   840 => x"1ee2d3c3",
   841 => x"fefe4974",
   842 => x"8ee887c8",
   843 => x"1e87d1fa",
   844 => x"c287d3fa",
   845 => x"c71ec11e",
   846 => x"d2fffe49",
   847 => x"c11ec287",
   848 => x"fe49c71e",
   849 => x"c087c8ff",
   850 => x"268ef048",
   851 => x"f2ebf44f",
   852 => x"040605f5",
   853 => x"830b030c",
   854 => x"fc00660a",
   855 => x"da005a00",
   856 => x"94800000",
   857 => x"78800508",
   858 => x"01800200",
   859 => x"09800300",
   860 => x"00800400",
   861 => x"91800100",
   862 => x"04002608",
   863 => x"00001d00",
   864 => x"00001c00",
   865 => x"0c002500",
   866 => x"00001a00",
   867 => x"00001b00",
   868 => x"00002400",
   869 => x"00011200",
   870 => x"03002e00",
   871 => x"00002d00",
   872 => x"00002300",
   873 => x"0b003600",
   874 => x"00002100",
   875 => x"00002b00",
   876 => x"00002c00",
   877 => x"00002200",
   878 => x"6c003d00",
   879 => x"00003500",
   880 => x"00003400",
   881 => x"75003e00",
   882 => x"00003200",
   883 => x"00003300",
   884 => x"6b003c00",
   885 => x"00002a00",
   886 => x"01004600",
   887 => x"73004300",
   888 => x"69003b00",
   889 => x"09004500",
   890 => x"70003a00",
   891 => x"72004200",
   892 => x"74004400",
   893 => x"00003100",
   894 => x"00005500",
   895 => x"7c004d00",
   896 => x"7a004b00",
   897 => x"00007b00",
   898 => x"71004900",
   899 => x"84004c00",
   900 => x"77005400",
   901 => x"00004100",
   902 => x"00006100",
   903 => x"7c005b00",
   904 => x"00005200",
   905 => x"0000f100",
   906 => x"00025900",
   907 => x"5d000e00",
   908 => x"00005d00",
   909 => x"79004a00",
   910 => x"05001600",
   911 => x"07007600",
   912 => x"0d000d00",
   913 => x"06001e00",
   914 => x"00002900",
   915 => x"00009100",
   916 => x"00001500",
   917 => x"00400000",
   918 => x"00008000",
   919 => x"00008000",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
