library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom1 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"f4d3c387",
    12 => x"86c0c64e",
    13 => x"49f4d3c3",
    14 => x"48e0f9c2",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087ede2",
    19 => x"1e87fc98",
    20 => x"1e731e72",
    21 => x"02114812",
    22 => x"c34b87ca",
    23 => x"739b98df",
    24 => x"87f00288",
    25 => x"4a264b26",
    26 => x"731e4f26",
    27 => x"c11e721e",
    28 => x"87ca048b",
    29 => x"02114812",
    30 => x"028887c4",
    31 => x"4a2687f1",
    32 => x"4f264b26",
    33 => x"731e741e",
    34 => x"c11e721e",
    35 => x"87d0048b",
    36 => x"02114812",
    37 => x"c34c87ca",
    38 => x"749c98df",
    39 => x"87eb0288",
    40 => x"4b264a26",
    41 => x"4f264c26",
    42 => x"8148731e",
    43 => x"c502a973",
    44 => x"05531287",
    45 => x"4f2687f6",
    46 => x"4a66c41e",
    47 => x"51124871",
    48 => x"2687fb05",
    49 => x"1e731e4f",
    50 => x"c0029a72",
    51 => x"48c087e7",
    52 => x"a9724bc1",
    53 => x"7287d106",
    54 => x"87c90682",
    55 => x"a9728373",
    56 => x"c387f401",
    57 => x"3ab2c187",
    58 => x"8903a972",
    59 => x"c1078073",
    60 => x"f3052b2a",
    61 => x"264b2687",
    62 => x"1e751e4f",
    63 => x"b7714dc4",
    64 => x"b9ff04a1",
    65 => x"bdc381c1",
    66 => x"a2b77207",
    67 => x"c1baff04",
    68 => x"07bdc182",
    69 => x"c187eefe",
    70 => x"b8ff042d",
    71 => x"2d0780c1",
    72 => x"c1b9ff04",
    73 => x"4d260781",
    74 => x"111e4f26",
    75 => x"08d4ff48",
    76 => x"4866c478",
    77 => x"a6c888c1",
    78 => x"05987058",
    79 => x"4f2687ed",
    80 => x"48d4ff1e",
    81 => x"6878ffc3",
    82 => x"4866c451",
    83 => x"a6c888c1",
    84 => x"05987058",
    85 => x"4f2687eb",
    86 => x"ff1e731e",
    87 => x"ffc34bd4",
    88 => x"c34a6b7b",
    89 => x"496b7bff",
    90 => x"b17232c8",
    91 => x"6b7bffc3",
    92 => x"7131c84a",
    93 => x"7bffc3b2",
    94 => x"32c8496b",
    95 => x"4871b172",
    96 => x"4d2687c4",
    97 => x"4b264c26",
    98 => x"5e0e4f26",
    99 => x"0e5d5c5b",
   100 => x"d4ff4a71",
   101 => x"c349724c",
   102 => x"7c7199ff",
   103 => x"bfe0f9c2",
   104 => x"d087c805",
   105 => x"30c94866",
   106 => x"d058a6d4",
   107 => x"29d84966",
   108 => x"7199ffc3",
   109 => x"4966d07c",
   110 => x"ffc329d0",
   111 => x"d07c7199",
   112 => x"29c84966",
   113 => x"7199ffc3",
   114 => x"4966d07c",
   115 => x"7199ffc3",
   116 => x"d049727c",
   117 => x"99ffc329",
   118 => x"4b6c7c71",
   119 => x"4dfff0c9",
   120 => x"05abffc3",
   121 => x"ffc387d0",
   122 => x"c14b6c7c",
   123 => x"87c6028d",
   124 => x"02abffc3",
   125 => x"487387f0",
   126 => x"1e87c7fe",
   127 => x"d4ff49c0",
   128 => x"78ffc348",
   129 => x"c8c381c1",
   130 => x"f104a9b7",
   131 => x"1e4f2687",
   132 => x"87e71e73",
   133 => x"4bdff8c4",
   134 => x"ffc01ec0",
   135 => x"49f7c1f0",
   136 => x"c487e7fd",
   137 => x"05a8c186",
   138 => x"ff87eac0",
   139 => x"ffc348d4",
   140 => x"c0c0c178",
   141 => x"1ec0c0c0",
   142 => x"c1f0e1c0",
   143 => x"c9fd49e9",
   144 => x"7086c487",
   145 => x"87ca0598",
   146 => x"c348d4ff",
   147 => x"48c178ff",
   148 => x"e6fe87cb",
   149 => x"058bc187",
   150 => x"c087fdfe",
   151 => x"87e6fc48",
   152 => x"ff1e731e",
   153 => x"ffc348d4",
   154 => x"c04bd378",
   155 => x"f0ffc01e",
   156 => x"fc49c1c1",
   157 => x"86c487d4",
   158 => x"ca059870",
   159 => x"48d4ff87",
   160 => x"c178ffc3",
   161 => x"fd87cb48",
   162 => x"8bc187f1",
   163 => x"87dbff05",
   164 => x"f1fb48c0",
   165 => x"5b5e0e87",
   166 => x"d4ff0e5c",
   167 => x"87dbfd4c",
   168 => x"c01eeac6",
   169 => x"c8c1f0e1",
   170 => x"87defb49",
   171 => x"a8c186c4",
   172 => x"fe87c802",
   173 => x"48c087ea",
   174 => x"fa87e2c1",
   175 => x"497087da",
   176 => x"99ffffcf",
   177 => x"02a9eac6",
   178 => x"d3fe87c8",
   179 => x"c148c087",
   180 => x"ffc387cb",
   181 => x"4bf1c07c",
   182 => x"7087f4fc",
   183 => x"ebc00298",
   184 => x"c01ec087",
   185 => x"fac1f0ff",
   186 => x"87defa49",
   187 => x"987086c4",
   188 => x"c387d905",
   189 => x"496c7cff",
   190 => x"7c7cffc3",
   191 => x"c0c17c7c",
   192 => x"87c40299",
   193 => x"87d548c1",
   194 => x"87d148c0",
   195 => x"c405abc2",
   196 => x"c848c087",
   197 => x"058bc187",
   198 => x"c087fdfe",
   199 => x"87e4f948",
   200 => x"c21e731e",
   201 => x"c148e0f9",
   202 => x"ff4bc778",
   203 => x"78c248d0",
   204 => x"ff87c8fb",
   205 => x"78c348d0",
   206 => x"e5c01ec0",
   207 => x"49c0c1d0",
   208 => x"c487c7f9",
   209 => x"05a8c186",
   210 => x"c24b87c1",
   211 => x"87c505ab",
   212 => x"f9c048c0",
   213 => x"058bc187",
   214 => x"fc87d0ff",
   215 => x"f9c287f7",
   216 => x"987058e4",
   217 => x"c187cd05",
   218 => x"f0ffc01e",
   219 => x"f849d0c1",
   220 => x"86c487d8",
   221 => x"c348d4ff",
   222 => x"e0c478ff",
   223 => x"e8f9c287",
   224 => x"48d0ff58",
   225 => x"d4ff78c2",
   226 => x"78ffc348",
   227 => x"f5f748c1",
   228 => x"5b5e0e87",
   229 => x"710e5d5c",
   230 => x"4dffc34a",
   231 => x"754cd4ff",
   232 => x"48d0ff7c",
   233 => x"7578c3c4",
   234 => x"c01e727c",
   235 => x"d8c1f0ff",
   236 => x"87d6f749",
   237 => x"987086c4",
   238 => x"c087c502",
   239 => x"87f0c048",
   240 => x"fec37c75",
   241 => x"1ec0c87c",
   242 => x"f54966d4",
   243 => x"86c487dc",
   244 => x"7c757c75",
   245 => x"dad87c75",
   246 => x"7c754be0",
   247 => x"0599496c",
   248 => x"8bc187c5",
   249 => x"7587f305",
   250 => x"48d0ff7c",
   251 => x"48c178c2",
   252 => x"1e87cff6",
   253 => x"ff4ad4ff",
   254 => x"d1c448d0",
   255 => x"7affc378",
   256 => x"f80589c1",
   257 => x"1e4f2687",
   258 => x"4b711e73",
   259 => x"dfcdeec5",
   260 => x"48d4ff4a",
   261 => x"6878ffc3",
   262 => x"a8fec348",
   263 => x"c187c502",
   264 => x"87ed058a",
   265 => x"c5059a72",
   266 => x"c048c087",
   267 => x"9b7387ea",
   268 => x"c887cc02",
   269 => x"49731e66",
   270 => x"c487c5f4",
   271 => x"c887c686",
   272 => x"eefe4966",
   273 => x"48d4ff87",
   274 => x"7878ffc3",
   275 => x"c5059b73",
   276 => x"48d0ff87",
   277 => x"48c178d0",
   278 => x"1e87ebf4",
   279 => x"4a711e73",
   280 => x"d4ff4bc0",
   281 => x"78ffc348",
   282 => x"c448d0ff",
   283 => x"d4ff78c3",
   284 => x"78ffc348",
   285 => x"ffc01e72",
   286 => x"49d1c1f0",
   287 => x"c487cbf4",
   288 => x"05987086",
   289 => x"c0c887cd",
   290 => x"4966cc1e",
   291 => x"c487f8fd",
   292 => x"ff4b7086",
   293 => x"78c248d0",
   294 => x"e9f34873",
   295 => x"5b5e0e87",
   296 => x"c00e5d5c",
   297 => x"f0ffc01e",
   298 => x"f349c9c1",
   299 => x"1ed287dc",
   300 => x"49e8f9c2",
   301 => x"c887d0fd",
   302 => x"c14cc086",
   303 => x"acb7d284",
   304 => x"c287f804",
   305 => x"bf97e8f9",
   306 => x"99c0c349",
   307 => x"05a9c0c1",
   308 => x"c287e7c0",
   309 => x"bf97eff9",
   310 => x"c231d049",
   311 => x"bf97f0f9",
   312 => x"7232c84a",
   313 => x"f1f9c2b1",
   314 => x"b14abf97",
   315 => x"ffcf4c71",
   316 => x"c19cffff",
   317 => x"c134ca84",
   318 => x"f9c287e7",
   319 => x"49bf97f1",
   320 => x"99c631c1",
   321 => x"97f2f9c2",
   322 => x"b7c74abf",
   323 => x"c2b1722a",
   324 => x"bf97edf9",
   325 => x"9dcf4d4a",
   326 => x"97eef9c2",
   327 => x"9ac34abf",
   328 => x"f9c232ca",
   329 => x"4bbf97ef",
   330 => x"b27333c2",
   331 => x"97f0f9c2",
   332 => x"c0c34bbf",
   333 => x"2bb7c69b",
   334 => x"81c2b273",
   335 => x"307148c1",
   336 => x"48c14970",
   337 => x"4d703075",
   338 => x"84c14c72",
   339 => x"c0c89471",
   340 => x"cc06adb7",
   341 => x"b734c187",
   342 => x"b7c0c82d",
   343 => x"f4ff01ad",
   344 => x"f0487487",
   345 => x"5e0e87dc",
   346 => x"0e5d5c5b",
   347 => x"c2c386f8",
   348 => x"78c048ce",
   349 => x"1ec6fac2",
   350 => x"defb49c0",
   351 => x"7086c487",
   352 => x"87c50598",
   353 => x"cec948c0",
   354 => x"c14dc087",
   355 => x"f8f9c07e",
   356 => x"fac249bf",
   357 => x"c8714afc",
   358 => x"87ceeb4b",
   359 => x"c2059870",
   360 => x"c07ec087",
   361 => x"49bff4f9",
   362 => x"4ad8fbc2",
   363 => x"ea4bc871",
   364 => x"987087f8",
   365 => x"c087c205",
   366 => x"c0026e7e",
   367 => x"c1c387fd",
   368 => x"c34dbfcc",
   369 => x"bf9fc4c2",
   370 => x"d6c5487e",
   371 => x"c705a8ea",
   372 => x"ccc1c387",
   373 => x"87ce4dbf",
   374 => x"e9ca486e",
   375 => x"c502a8d5",
   376 => x"c748c087",
   377 => x"fac287f1",
   378 => x"49751ec6",
   379 => x"c487ecf9",
   380 => x"05987086",
   381 => x"48c087c5",
   382 => x"c087dcc7",
   383 => x"49bff4f9",
   384 => x"4ad8fbc2",
   385 => x"e94bc871",
   386 => x"987087e0",
   387 => x"c387c805",
   388 => x"c148cec2",
   389 => x"c087da78",
   390 => x"49bff8f9",
   391 => x"4afcfac2",
   392 => x"e94bc871",
   393 => x"987087c4",
   394 => x"87c5c002",
   395 => x"e6c648c0",
   396 => x"c4c2c387",
   397 => x"c149bf97",
   398 => x"c005a9d5",
   399 => x"c2c387cd",
   400 => x"49bf97c5",
   401 => x"02a9eac2",
   402 => x"c087c5c0",
   403 => x"87c7c648",
   404 => x"97c6fac2",
   405 => x"c3487ebf",
   406 => x"c002a8e9",
   407 => x"486e87ce",
   408 => x"02a8ebc3",
   409 => x"c087c5c0",
   410 => x"87ebc548",
   411 => x"97d1fac2",
   412 => x"059949bf",
   413 => x"c287ccc0",
   414 => x"bf97d2fa",
   415 => x"02a9c249",
   416 => x"c087c5c0",
   417 => x"87cfc548",
   418 => x"97d3fac2",
   419 => x"c2c348bf",
   420 => x"4c7058ca",
   421 => x"c388c148",
   422 => x"c258cec2",
   423 => x"bf97d4fa",
   424 => x"c2817549",
   425 => x"bf97d5fa",
   426 => x"7232c84a",
   427 => x"c6c37ea1",
   428 => x"786e48db",
   429 => x"97d6fac2",
   430 => x"a6c848bf",
   431 => x"cec2c358",
   432 => x"d4c202bf",
   433 => x"f4f9c087",
   434 => x"fbc249bf",
   435 => x"c8714ad8",
   436 => x"87d6e64b",
   437 => x"c0029870",
   438 => x"48c087c5",
   439 => x"c387f8c3",
   440 => x"4cbfc6c2",
   441 => x"5cefc6c3",
   442 => x"97ebfac2",
   443 => x"31c849bf",
   444 => x"97eafac2",
   445 => x"49a14abf",
   446 => x"97ecfac2",
   447 => x"32d04abf",
   448 => x"c249a172",
   449 => x"bf97edfa",
   450 => x"7232d84a",
   451 => x"66c449a1",
   452 => x"dbc6c391",
   453 => x"c6c381bf",
   454 => x"fac259e3",
   455 => x"4abf97f3",
   456 => x"fac232c8",
   457 => x"4bbf97f2",
   458 => x"fac24aa2",
   459 => x"4bbf97f4",
   460 => x"a27333d0",
   461 => x"f5fac24a",
   462 => x"cf4bbf97",
   463 => x"7333d89b",
   464 => x"c6c34aa2",
   465 => x"c6c35ae7",
   466 => x"c24abfe3",
   467 => x"c392748a",
   468 => x"7248e7c6",
   469 => x"cac178a1",
   470 => x"d8fac287",
   471 => x"c849bf97",
   472 => x"d7fac231",
   473 => x"a14abf97",
   474 => x"d6c2c349",
   475 => x"d2c2c359",
   476 => x"31c549bf",
   477 => x"c981ffc7",
   478 => x"efc6c329",
   479 => x"ddfac259",
   480 => x"c84abf97",
   481 => x"dcfac232",
   482 => x"a24bbf97",
   483 => x"9266c44a",
   484 => x"c6c3826e",
   485 => x"c6c35aeb",
   486 => x"78c048e3",
   487 => x"48dfc6c3",
   488 => x"c378a172",
   489 => x"c348efc6",
   490 => x"78bfe3c6",
   491 => x"48f3c6c3",
   492 => x"bfe7c6c3",
   493 => x"cec2c378",
   494 => x"c9c002bf",
   495 => x"c4487487",
   496 => x"c07e7030",
   497 => x"c6c387c9",
   498 => x"c448bfeb",
   499 => x"c37e7030",
   500 => x"6e48d2c2",
   501 => x"f848c178",
   502 => x"264d268e",
   503 => x"264b264c",
   504 => x"5b5e0e4f",
   505 => x"710e5d5c",
   506 => x"cec2c34a",
   507 => x"87cb02bf",
   508 => x"2bc74b72",
   509 => x"ffc14c72",
   510 => x"7287c99c",
   511 => x"722bc84b",
   512 => x"9cffc34c",
   513 => x"bfdbc6c3",
   514 => x"f0f9c083",
   515 => x"d902abbf",
   516 => x"f4f9c087",
   517 => x"c6fac25b",
   518 => x"f049731e",
   519 => x"86c487fd",
   520 => x"c5059870",
   521 => x"c048c087",
   522 => x"c2c387e6",
   523 => x"d202bfce",
   524 => x"c4497487",
   525 => x"c6fac291",
   526 => x"cf4d6981",
   527 => x"ffffffff",
   528 => x"7487cb9d",
   529 => x"c291c249",
   530 => x"9f81c6fa",
   531 => x"48754d69",
   532 => x"0e87c6fe",
   533 => x"5d5c5b5e",
   534 => x"4d711e0e",
   535 => x"49c11ec0",
   536 => x"c487f5d0",
   537 => x"9c4c7086",
   538 => x"87c2c102",
   539 => x"4ad6c2c3",
   540 => x"dfff4975",
   541 => x"987087d9",
   542 => x"87f2c002",
   543 => x"49754a74",
   544 => x"dfff4bcb",
   545 => x"987087fe",
   546 => x"87e2c002",
   547 => x"9c741ec0",
   548 => x"c487c702",
   549 => x"78c048a6",
   550 => x"a6c487c5",
   551 => x"c478c148",
   552 => x"f3cf4966",
   553 => x"7086c487",
   554 => x"fe059c4c",
   555 => x"487487fe",
   556 => x"87e5fc26",
   557 => x"5c5b5e0e",
   558 => x"86f80e5d",
   559 => x"059b4b71",
   560 => x"48c087c5",
   561 => x"c887d4c2",
   562 => x"7dc04da3",
   563 => x"c70266d8",
   564 => x"9766d887",
   565 => x"87c505bf",
   566 => x"fec148c0",
   567 => x"4966d887",
   568 => x"7087f0fd",
   569 => x"c1026e7e",
   570 => x"496e87ef",
   571 => x"7d6981dc",
   572 => x"81da496e",
   573 => x"9f4ca3c4",
   574 => x"c2c37c69",
   575 => x"d002bfce",
   576 => x"d4496e87",
   577 => x"49699f81",
   578 => x"ffffc04a",
   579 => x"c232d09a",
   580 => x"724ac087",
   581 => x"806c4849",
   582 => x"7bc07c70",
   583 => x"6c49a3cc",
   584 => x"49a3d079",
   585 => x"a6c479c0",
   586 => x"d478c048",
   587 => x"66c44aa3",
   588 => x"7291c849",
   589 => x"41c049a1",
   590 => x"66c4796c",
   591 => x"c880c148",
   592 => x"b7d058a6",
   593 => x"e2ff04a8",
   594 => x"c94a6d87",
   595 => x"c22ac72a",
   596 => x"7249a3d4",
   597 => x"c2486e79",
   598 => x"f848c087",
   599 => x"87f9f98e",
   600 => x"5c5b5e0e",
   601 => x"4c710e5d",
   602 => x"48f0f9c0",
   603 => x"9c7478ff",
   604 => x"87cac102",
   605 => x"6949a4c8",
   606 => x"87c2c102",
   607 => x"6c4a66d0",
   608 => x"a6d48249",
   609 => x"4d66d05a",
   610 => x"cac2c3b9",
   611 => x"baff4abf",
   612 => x"99719972",
   613 => x"87e4c002",
   614 => x"6b4ba4c4",
   615 => x"87c1f949",
   616 => x"c2c37b70",
   617 => x"6c49bfc6",
   618 => x"757c7181",
   619 => x"cac2c3b9",
   620 => x"baff4abf",
   621 => x"99719972",
   622 => x"87dcff05",
   623 => x"d8f87c75",
   624 => x"1e731e87",
   625 => x"029b4b71",
   626 => x"a3c887c7",
   627 => x"c5056949",
   628 => x"c048c087",
   629 => x"c6c387eb",
   630 => x"c44abfdf",
   631 => x"496949a3",
   632 => x"c2c389c2",
   633 => x"7191bfc6",
   634 => x"c2c34aa2",
   635 => x"6b49bfca",
   636 => x"4aa27199",
   637 => x"721e66c8",
   638 => x"87dfe949",
   639 => x"497086c4",
   640 => x"87d9f748",
   641 => x"711e731e",
   642 => x"c7029b4b",
   643 => x"49a3c887",
   644 => x"87c50569",
   645 => x"ebc048c0",
   646 => x"dfc6c387",
   647 => x"a3c44abf",
   648 => x"c2496949",
   649 => x"c6c2c389",
   650 => x"a27191bf",
   651 => x"cac2c34a",
   652 => x"996b49bf",
   653 => x"c84aa271",
   654 => x"49721e66",
   655 => x"c487d2e5",
   656 => x"48497086",
   657 => x"0e87d6f6",
   658 => x"5d5c5b5e",
   659 => x"7186f80e",
   660 => x"48a6c44b",
   661 => x"a3c878ff",
   662 => x"c04d6949",
   663 => x"4aa3d44c",
   664 => x"91c84974",
   665 => x"6949a172",
   666 => x"4866d849",
   667 => x"7e708871",
   668 => x"01a966d8",
   669 => x"ad6e87ca",
   670 => x"c887c506",
   671 => x"4d6e5ca6",
   672 => x"b7d084c1",
   673 => x"d4ff04ac",
   674 => x"4866c487",
   675 => x"c8f58ef8",
   676 => x"5b5e0e87",
   677 => x"ec0e5d5c",
   678 => x"59a6c886",
   679 => x"c148a6c8",
   680 => x"ffffffff",
   681 => x"80c478ff",
   682 => x"4dc078ff",
   683 => x"66c44cc0",
   684 => x"7483d44b",
   685 => x"7391c849",
   686 => x"4a7549a1",
   687 => x"a27392c8",
   688 => x"6e49697e",
   689 => x"a6d489bf",
   690 => x"05ad7459",
   691 => x"a6d087c6",
   692 => x"78bf6e48",
   693 => x"c04866d0",
   694 => x"cf04a8b7",
   695 => x"4966d087",
   696 => x"03a966c8",
   697 => x"a6d087c6",
   698 => x"59a6cc5c",
   699 => x"b7d084c1",
   700 => x"f9fe04ac",
   701 => x"d085c187",
   702 => x"fe04adb7",
   703 => x"66cc87ee",
   704 => x"f38eec48",
   705 => x"5e0e87d3",
   706 => x"0e5d5c5b",
   707 => x"4b7186f0",
   708 => x"4c66e0c0",
   709 => x"9b732cc9",
   710 => x"87e1c302",
   711 => x"6949a3c8",
   712 => x"87d9c302",
   713 => x"c049a3d0",
   714 => x"6b7966e0",
   715 => x"c302ac7e",
   716 => x"c2c387cb",
   717 => x"ff49bfca",
   718 => x"744a71b9",
   719 => x"6e48719a",
   720 => x"58a6cc98",
   721 => x"c44da3c4",
   722 => x"786d48a6",
   723 => x"05aa66c8",
   724 => x"7b7487c5",
   725 => x"7287d1c2",
   726 => x"fb49731e",
   727 => x"86c487e9",
   728 => x"c0487e70",
   729 => x"d004a8b7",
   730 => x"4aa3d487",
   731 => x"91c8496e",
   732 => x"2149a172",
   733 => x"c77d697b",
   734 => x"cc7bc087",
   735 => x"7d6949a3",
   736 => x"731e66c8",
   737 => x"87fffa49",
   738 => x"7e7086c4",
   739 => x"49a3d4c2",
   740 => x"6948a6cc",
   741 => x"4866c878",
   742 => x"06a866cc",
   743 => x"486e87c9",
   744 => x"04a8b7c0",
   745 => x"6e87e0c0",
   746 => x"a8b7c048",
   747 => x"87ecc004",
   748 => x"6e4aa3d4",
   749 => x"7291c849",
   750 => x"66c849a1",
   751 => x"70886948",
   752 => x"a966cc49",
   753 => x"7387d506",
   754 => x"87c5fb49",
   755 => x"a3d44970",
   756 => x"7291c84a",
   757 => x"66c849a1",
   758 => x"7966c441",
   759 => x"49748c6b",
   760 => x"f549731e",
   761 => x"86c487fa",
   762 => x"4966e0c0",
   763 => x"0299ffc7",
   764 => x"fac287cb",
   765 => x"49731ec6",
   766 => x"c487c6f7",
   767 => x"ef8ef086",
   768 => x"731e87d7",
   769 => x"9b4b711e",
   770 => x"87e4c002",
   771 => x"5bf3c6c3",
   772 => x"8ac24a73",
   773 => x"bfc6c2c3",
   774 => x"c6c39249",
   775 => x"7248bfdf",
   776 => x"f7c6c380",
   777 => x"c4487158",
   778 => x"d6c2c330",
   779 => x"87edc058",
   780 => x"48efc6c3",
   781 => x"bfe3c6c3",
   782 => x"f3c6c378",
   783 => x"e7c6c348",
   784 => x"c2c378bf",
   785 => x"c902bfce",
   786 => x"c6c2c387",
   787 => x"31c449bf",
   788 => x"c6c387c7",
   789 => x"c449bfeb",
   790 => x"d6c2c331",
   791 => x"87fded59",
   792 => x"5c5b5e0e",
   793 => x"c04a710e",
   794 => x"029a724b",
   795 => x"da87e1c0",
   796 => x"699f49a2",
   797 => x"cec2c34b",
   798 => x"87cf02bf",
   799 => x"9f49a2d4",
   800 => x"c04c4969",
   801 => x"d09cffff",
   802 => x"c087c234",
   803 => x"b349744c",
   804 => x"edfd4973",
   805 => x"87c3ed87",
   806 => x"5c5b5e0e",
   807 => x"86f40e5d",
   808 => x"7ec04a71",
   809 => x"d8029a72",
   810 => x"c2fac287",
   811 => x"c278c048",
   812 => x"c348faf9",
   813 => x"78bff3c6",
   814 => x"48fef9c2",
   815 => x"bfefc6c3",
   816 => x"e3c2c378",
   817 => x"c350c048",
   818 => x"49bfd2c2",
   819 => x"bfc2fac2",
   820 => x"03aa714a",
   821 => x"7287c0c4",
   822 => x"0599cf49",
   823 => x"c287e1c0",
   824 => x"c21ec6fa",
   825 => x"49bffaf9",
   826 => x"48faf9c2",
   827 => x"7178a1c1",
   828 => x"87e7ddff",
   829 => x"f9c086c4",
   830 => x"fac248ec",
   831 => x"87cc78c6",
   832 => x"bfecf9c0",
   833 => x"80e0c048",
   834 => x"58f0f9c0",
   835 => x"bfc2fac2",
   836 => x"c280c148",
   837 => x"2758c6fa",
   838 => x"00000e6c",
   839 => x"4dbf97bf",
   840 => x"e2c2029d",
   841 => x"ade5c387",
   842 => x"87dbc202",
   843 => x"bfecf9c0",
   844 => x"49a3cb4b",
   845 => x"accf4c11",
   846 => x"87d2c105",
   847 => x"99df4975",
   848 => x"91cd89c1",
   849 => x"81d6c2c3",
   850 => x"124aa3c1",
   851 => x"4aa3c351",
   852 => x"a3c55112",
   853 => x"c751124a",
   854 => x"51124aa3",
   855 => x"124aa3c9",
   856 => x"4aa3ce51",
   857 => x"a3d05112",
   858 => x"d251124a",
   859 => x"51124aa3",
   860 => x"124aa3d4",
   861 => x"4aa3d651",
   862 => x"a3d85112",
   863 => x"dc51124a",
   864 => x"51124aa3",
   865 => x"124aa3de",
   866 => x"c07ec151",
   867 => x"497487f9",
   868 => x"c00599c8",
   869 => x"497487ea",
   870 => x"d00599d0",
   871 => x"0266dc87",
   872 => x"7387cac0",
   873 => x"0f66dc49",
   874 => x"d3029870",
   875 => x"c0056e87",
   876 => x"c2c387c6",
   877 => x"50c048d6",
   878 => x"bfecf9c0",
   879 => x"87e7c248",
   880 => x"48e3c2c3",
   881 => x"c37e50c0",
   882 => x"49bfd2c2",
   883 => x"bfc2fac2",
   884 => x"04aa714a",
   885 => x"c387c0fc",
   886 => x"05bff3c6",
   887 => x"c387c8c0",
   888 => x"02bfcec2",
   889 => x"c087fec1",
   890 => x"ff48f0f9",
   891 => x"fef9c278",
   892 => x"ece749bf",
   893 => x"c2497087",
   894 => x"c459c2fa",
   895 => x"f9c248a6",
   896 => x"c378bffe",
   897 => x"02bfcec2",
   898 => x"c487d8c0",
   899 => x"ffcf4966",
   900 => x"99f8ffff",
   901 => x"c5c002a9",
   902 => x"c04dc087",
   903 => x"4dc187e1",
   904 => x"c487dcc0",
   905 => x"ffcf4966",
   906 => x"02a999f8",
   907 => x"c887c8c0",
   908 => x"78c048a6",
   909 => x"c887c5c0",
   910 => x"78c148a6",
   911 => x"754d66c8",
   912 => x"e0c0059d",
   913 => x"4966c487",
   914 => x"c2c389c2",
   915 => x"914abfc6",
   916 => x"bfdfc6c3",
   917 => x"faf9c24a",
   918 => x"78a17248",
   919 => x"48c2fac2",
   920 => x"e2f978c0",
   921 => x"f448c087",
   922 => x"87ede58e",
   923 => x"00000000",
   924 => x"ffffffff",
   925 => x"00000e7c",
   926 => x"00000e85",
   927 => x"33544146",
   928 => x"20202032",
   929 => x"54414600",
   930 => x"20203631",
   931 => x"ff1e0020",
   932 => x"ffc348d4",
   933 => x"26486878",
   934 => x"d4ff1e4f",
   935 => x"78ffc348",
   936 => x"c848d0ff",
   937 => x"d4ff78e1",
   938 => x"c378d448",
   939 => x"ff48f7c6",
   940 => x"2650bfd4",
   941 => x"d0ff1e4f",
   942 => x"78e0c048",
   943 => x"ff1e4f26",
   944 => x"497087cc",
   945 => x"87c60299",
   946 => x"05a9fbc0",
   947 => x"487187f1",
   948 => x"5e0e4f26",
   949 => x"710e5c5b",
   950 => x"fe4cc04b",
   951 => x"497087f0",
   952 => x"f9c00299",
   953 => x"a9ecc087",
   954 => x"87f2c002",
   955 => x"02a9fbc0",
   956 => x"cc87ebc0",
   957 => x"03acb766",
   958 => x"66d087c7",
   959 => x"7187c202",
   960 => x"02997153",
   961 => x"84c187c2",
   962 => x"7087c3fe",
   963 => x"cd029949",
   964 => x"a9ecc087",
   965 => x"c087c702",
   966 => x"ff05a9fb",
   967 => x"66d087d5",
   968 => x"c087c302",
   969 => x"ecc07b97",
   970 => x"87c405a9",
   971 => x"87c54a74",
   972 => x"0ac04a74",
   973 => x"c248728a",
   974 => x"264d2687",
   975 => x"264b264c",
   976 => x"c9fd1e4f",
   977 => x"c0497087",
   978 => x"04a9b7f0",
   979 => x"f9c087ca",
   980 => x"c301a9b7",
   981 => x"89f0c087",
   982 => x"a9b7c1c1",
   983 => x"c187ca04",
   984 => x"01a9b7da",
   985 => x"f7c087c3",
   986 => x"26487189",
   987 => x"5b5e0e4f",
   988 => x"4a710e5c",
   989 => x"724cd4ff",
   990 => x"87eac049",
   991 => x"029b4b70",
   992 => x"8bc187c2",
   993 => x"c848d0ff",
   994 => x"d5c178c5",
   995 => x"c649737c",
   996 => x"c5e2c231",
   997 => x"484abf97",
   998 => x"7c70b071",
   999 => x"c448d0ff",
  1000 => x"fe487378",
  1001 => x"5e0e87d5",
  1002 => x"0e5d5c5b",
  1003 => x"4c7186f8",
  1004 => x"e4fb7ec0",
  1005 => x"c14bc087",
  1006 => x"bf97d3c1",
  1007 => x"04a9c049",
  1008 => x"f9fb87cf",
  1009 => x"c183c187",
  1010 => x"bf97d3c1",
  1011 => x"f106ab49",
  1012 => x"d3c1c187",
  1013 => x"cf02bf97",
  1014 => x"87f2fa87",
  1015 => x"02994970",
  1016 => x"ecc087c6",
  1017 => x"87f105a9",
  1018 => x"e1fa4bc0",
  1019 => x"fa4d7087",
  1020 => x"a6c887dc",
  1021 => x"87d6fa58",
  1022 => x"83c14a70",
  1023 => x"9749a4c8",
  1024 => x"02ad4969",
  1025 => x"ffc087c7",
  1026 => x"e7c005ad",
  1027 => x"49a4c987",
  1028 => x"c4496997",
  1029 => x"c702a966",
  1030 => x"ffc04887",
  1031 => x"87d405a8",
  1032 => x"9749a4ca",
  1033 => x"02aa4969",
  1034 => x"ffc087c6",
  1035 => x"87c405aa",
  1036 => x"87d07ec1",
  1037 => x"02adecc0",
  1038 => x"fbc087c6",
  1039 => x"87c405ad",
  1040 => x"7ec14bc0",
  1041 => x"e1fe026e",
  1042 => x"87e9f987",
  1043 => x"8ef84873",
  1044 => x"0087e6fb",
  1045 => x"5c5b5e0e",
  1046 => x"711e0e5d",
  1047 => x"4d4cc04b",
  1048 => x"e8c004ab",
  1049 => x"e6fec087",
  1050 => x"029d751e",
  1051 => x"4ac087c4",
  1052 => x"4ac187c2",
  1053 => x"dff04972",
  1054 => x"7086c487",
  1055 => x"6e84c17e",
  1056 => x"7387c205",
  1057 => x"7385c14c",
  1058 => x"d8ff06ac",
  1059 => x"26486e87",
  1060 => x"4c264d26",
  1061 => x"4f264b26",
  1062 => x"5c5b5e0e",
  1063 => x"711e0e5d",
  1064 => x"91de494c",
  1065 => x"4dd1c7c3",
  1066 => x"6d978571",
  1067 => x"87ddc102",
  1068 => x"bffcc6c3",
  1069 => x"7282744a",
  1070 => x"87d8fe49",
  1071 => x"026e7e70",
  1072 => x"c387f3c0",
  1073 => x"6e4bc4c7",
  1074 => x"fe49cb4a",
  1075 => x"7487d9ff",
  1076 => x"c193cb4b",
  1077 => x"c483dce4",
  1078 => x"d1c4c183",
  1079 => x"c149747b",
  1080 => x"7587fec2",
  1081 => x"d0c7c37b",
  1082 => x"1e49bf97",
  1083 => x"49c4c7c3",
  1084 => x"87d3ddc1",
  1085 => x"497486c4",
  1086 => x"87e5c2c1",
  1087 => x"c4c149c0",
  1088 => x"c6c387c4",
  1089 => x"78c048f8",
  1090 => x"fadc49c1",
  1091 => x"fffd2687",
  1092 => x"616f4c87",
  1093 => x"676e6964",
  1094 => x"002e2e2e",
  1095 => x"5c5b5e0e",
  1096 => x"4a4b710e",
  1097 => x"bffcc6c3",
  1098 => x"fc497282",
  1099 => x"4c7087e6",
  1100 => x"87c4029c",
  1101 => x"87e8ec49",
  1102 => x"48fcc6c3",
  1103 => x"49c178c0",
  1104 => x"fd87c4dc",
  1105 => x"5e0e87cc",
  1106 => x"0e5d5c5b",
  1107 => x"fac286f4",
  1108 => x"4cc04dc6",
  1109 => x"c048a6c4",
  1110 => x"fcc6c378",
  1111 => x"a9c049bf",
  1112 => x"87c1c106",
  1113 => x"48c6fac2",
  1114 => x"f8c00298",
  1115 => x"e6fec087",
  1116 => x"0266c81e",
  1117 => x"a6c487c7",
  1118 => x"c578c048",
  1119 => x"48a6c487",
  1120 => x"66c478c1",
  1121 => x"87d0ec49",
  1122 => x"4d7086c4",
  1123 => x"66c484c1",
  1124 => x"c880c148",
  1125 => x"c6c358a6",
  1126 => x"ac49bffc",
  1127 => x"7587c603",
  1128 => x"c8ff059d",
  1129 => x"754cc087",
  1130 => x"e0c3029d",
  1131 => x"e6fec087",
  1132 => x"0266c81e",
  1133 => x"a6cc87c7",
  1134 => x"c578c048",
  1135 => x"48a6cc87",
  1136 => x"66cc78c1",
  1137 => x"87d0eb49",
  1138 => x"7e7086c4",
  1139 => x"e9c2026e",
  1140 => x"cb496e87",
  1141 => x"49699781",
  1142 => x"c10299d0",
  1143 => x"c4c187d6",
  1144 => x"49744adc",
  1145 => x"e4c191cb",
  1146 => x"797281dc",
  1147 => x"ffc381c8",
  1148 => x"de497451",
  1149 => x"d1c7c391",
  1150 => x"c285714d",
  1151 => x"c17d97c1",
  1152 => x"e0c049a5",
  1153 => x"d6c2c351",
  1154 => x"d202bf97",
  1155 => x"c284c187",
  1156 => x"c2c34ba5",
  1157 => x"49db4ad6",
  1158 => x"87ccfafe",
  1159 => x"cd87dbc1",
  1160 => x"51c049a5",
  1161 => x"a5c284c1",
  1162 => x"cb4a6e4b",
  1163 => x"f7f9fe49",
  1164 => x"87c6c187",
  1165 => x"4ad8c2c1",
  1166 => x"91cb4974",
  1167 => x"81dce4c1",
  1168 => x"c2c37972",
  1169 => x"02bf97d6",
  1170 => x"497487d8",
  1171 => x"84c191de",
  1172 => x"4bd1c7c3",
  1173 => x"c2c38371",
  1174 => x"49dd4ad6",
  1175 => x"87c8f9fe",
  1176 => x"4b7487d8",
  1177 => x"c7c393de",
  1178 => x"a3cb83d1",
  1179 => x"c151c049",
  1180 => x"4a6e7384",
  1181 => x"f8fe49cb",
  1182 => x"66c487ee",
  1183 => x"c880c148",
  1184 => x"acc758a6",
  1185 => x"87c5c003",
  1186 => x"e0fc056e",
  1187 => x"f4487487",
  1188 => x"87fcf78e",
  1189 => x"711e731e",
  1190 => x"91cb494b",
  1191 => x"81dce4c1",
  1192 => x"c24aa1c8",
  1193 => x"1248c5e2",
  1194 => x"4aa1c950",
  1195 => x"48d3c1c1",
  1196 => x"81ca5012",
  1197 => x"48d0c7c3",
  1198 => x"c7c35011",
  1199 => x"49bf97d0",
  1200 => x"c149c01e",
  1201 => x"c387c0d6",
  1202 => x"de48f8c6",
  1203 => x"d549c178",
  1204 => x"f62687f5",
  1205 => x"711e87fe",
  1206 => x"91cb494a",
  1207 => x"81dce4c1",
  1208 => x"481181c8",
  1209 => x"58fcc6c3",
  1210 => x"48fcc6c3",
  1211 => x"49c178c0",
  1212 => x"2687d4d5",
  1213 => x"49c01e4f",
  1214 => x"87cafcc0",
  1215 => x"711e4f26",
  1216 => x"87d20299",
  1217 => x"48f1e5c1",
  1218 => x"80f750c0",
  1219 => x"40d6cbc1",
  1220 => x"78d5e4c1",
  1221 => x"e5c187ce",
  1222 => x"e4c148ed",
  1223 => x"80fc78ce",
  1224 => x"78f5cbc1",
  1225 => x"5e0e4f26",
  1226 => x"710e5c5b",
  1227 => x"92cb4a4c",
  1228 => x"82dce4c1",
  1229 => x"c949a2c8",
  1230 => x"6b974ba2",
  1231 => x"69971e4b",
  1232 => x"82ca1e49",
  1233 => x"e7c04912",
  1234 => x"49c087c5",
  1235 => x"7487f8d3",
  1236 => x"ccf9c049",
  1237 => x"f48ef887",
  1238 => x"731e87f8",
  1239 => x"c64b711e",
  1240 => x"db024aa3",
  1241 => x"028ac187",
  1242 => x"028a87d6",
  1243 => x"8a87dac1",
  1244 => x"87fcc002",
  1245 => x"e1c0028a",
  1246 => x"cb028a87",
  1247 => x"87dbc187",
  1248 => x"d1fd49c7",
  1249 => x"87dec187",
  1250 => x"bffcc6c3",
  1251 => x"87cbc102",
  1252 => x"c388c148",
  1253 => x"c158c0c7",
  1254 => x"c7c387c1",
  1255 => x"c002bfc0",
  1256 => x"c6c387f9",
  1257 => x"c148bffc",
  1258 => x"c0c7c380",
  1259 => x"87ebc058",
  1260 => x"bffcc6c3",
  1261 => x"c389c649",
  1262 => x"c059c0c7",
  1263 => x"da03a9b7",
  1264 => x"fcc6c387",
  1265 => x"d278c048",
  1266 => x"c0c7c387",
  1267 => x"87cb02bf",
  1268 => x"bffcc6c3",
  1269 => x"c380c648",
  1270 => x"c058c0c7",
  1271 => x"87e7d149",
  1272 => x"f6c04973",
  1273 => x"ebf287fb",
  1274 => x"5b5e0e87",
  1275 => x"4c710e5c",
  1276 => x"741e66cc",
  1277 => x"c193cb4b",
  1278 => x"c483dce4",
  1279 => x"496a4aa3",
  1280 => x"87f4f2fe",
  1281 => x"7bd4cac1",
  1282 => x"d449a3c8",
  1283 => x"a3c95166",
  1284 => x"5166d849",
  1285 => x"dc49a3ca",
  1286 => x"f1265166",
  1287 => x"5e0e87f4",
  1288 => x"0e5d5c5b",
  1289 => x"d886d0ff",
  1290 => x"a6c459a6",
  1291 => x"c478c048",
  1292 => x"66c4c180",
  1293 => x"c180c478",
  1294 => x"c180c478",
  1295 => x"c0c7c378",
  1296 => x"c378c148",
  1297 => x"48bff8c6",
  1298 => x"cb05a8de",
  1299 => x"87f6f387",
  1300 => x"a6c84970",
  1301 => x"87f8ce59",
  1302 => x"e987fee8",
  1303 => x"ede887e0",
  1304 => x"c04c7087",
  1305 => x"c102acfb",
  1306 => x"66d487d0",
  1307 => x"87c2c105",
  1308 => x"c11e1ec0",
  1309 => x"ffe5c11e",
  1310 => x"fd49c01e",
  1311 => x"d0c187eb",
  1312 => x"82c44a66",
  1313 => x"81c7496a",
  1314 => x"1ec15174",
  1315 => x"496a1ed8",
  1316 => x"fde881c8",
  1317 => x"c186d887",
  1318 => x"c04866c4",
  1319 => x"87c701a8",
  1320 => x"c148a6c4",
  1321 => x"c187ce78",
  1322 => x"c14866c4",
  1323 => x"58a6cc88",
  1324 => x"c9e887c3",
  1325 => x"48a6cc87",
  1326 => x"9c7478c2",
  1327 => x"87cccd02",
  1328 => x"c14866c4",
  1329 => x"03a866c8",
  1330 => x"d887c1cd",
  1331 => x"78c048a6",
  1332 => x"7087fbe6",
  1333 => x"acd0c14c",
  1334 => x"87d6c205",
  1335 => x"e97e66d8",
  1336 => x"497087df",
  1337 => x"e659a6dc",
  1338 => x"4c7087e4",
  1339 => x"05acecc0",
  1340 => x"c487eac1",
  1341 => x"91cb4966",
  1342 => x"8166c0c1",
  1343 => x"6a4aa1c4",
  1344 => x"4aa1c84d",
  1345 => x"c15266d8",
  1346 => x"e679d6cb",
  1347 => x"4c7087c0",
  1348 => x"87d8029c",
  1349 => x"02acfbc0",
  1350 => x"557487d2",
  1351 => x"7087efe5",
  1352 => x"c7029c4c",
  1353 => x"acfbc087",
  1354 => x"87eeff05",
  1355 => x"c255e0c0",
  1356 => x"97c055c1",
  1357 => x"4966d47d",
  1358 => x"db05a96e",
  1359 => x"4866c487",
  1360 => x"04a866c8",
  1361 => x"66c487ca",
  1362 => x"c880c148",
  1363 => x"87c858a6",
  1364 => x"c14866c8",
  1365 => x"58a6cc88",
  1366 => x"7087f3e4",
  1367 => x"acd0c14c",
  1368 => x"d087c805",
  1369 => x"80c14866",
  1370 => x"c158a6d4",
  1371 => x"fd02acd0",
  1372 => x"a6dc87ea",
  1373 => x"7866d448",
  1374 => x"dc4866d8",
  1375 => x"c905a866",
  1376 => x"e0c087dc",
  1377 => x"f0c048a6",
  1378 => x"cc80c478",
  1379 => x"80c47866",
  1380 => x"747e78c0",
  1381 => x"88fbc048",
  1382 => x"58a6f0c0",
  1383 => x"c8029870",
  1384 => x"cb4887d7",
  1385 => x"a6f0c088",
  1386 => x"02987058",
  1387 => x"4887e9c0",
  1388 => x"f0c088c9",
  1389 => x"987058a6",
  1390 => x"87e1c302",
  1391 => x"c088c448",
  1392 => x"7058a6f0",
  1393 => x"87de0298",
  1394 => x"c088c148",
  1395 => x"7058a6f0",
  1396 => x"c8c30298",
  1397 => x"87dbc787",
  1398 => x"48a6e0c0",
  1399 => x"66cc78c0",
  1400 => x"d080c148",
  1401 => x"e5e258a6",
  1402 => x"c04c7087",
  1403 => x"d502acec",
  1404 => x"66e0c087",
  1405 => x"c087c602",
  1406 => x"c95ca6e4",
  1407 => x"c0487487",
  1408 => x"e8c088f0",
  1409 => x"ecc058a6",
  1410 => x"87cc02ac",
  1411 => x"7087ffe1",
  1412 => x"acecc04c",
  1413 => x"87f4ff05",
  1414 => x"1e66e0c0",
  1415 => x"1e4966d4",
  1416 => x"1e66ecc0",
  1417 => x"1effe5c1",
  1418 => x"f64966d4",
  1419 => x"1ec087fb",
  1420 => x"66dc1eca",
  1421 => x"c191cb49",
  1422 => x"d88166d8",
  1423 => x"a1c448a6",
  1424 => x"bf66d878",
  1425 => x"87cae249",
  1426 => x"b7c086d8",
  1427 => x"c7c106a8",
  1428 => x"de1ec187",
  1429 => x"bf66c81e",
  1430 => x"87f6e149",
  1431 => x"497086c8",
  1432 => x"8808c048",
  1433 => x"58a6e4c0",
  1434 => x"06a8b7c0",
  1435 => x"c087e9c0",
  1436 => x"dd4866e0",
  1437 => x"df03a8b7",
  1438 => x"49bf6e87",
  1439 => x"8166e0c0",
  1440 => x"6651e0c0",
  1441 => x"6e81c149",
  1442 => x"c1c281bf",
  1443 => x"66e0c051",
  1444 => x"6e81c249",
  1445 => x"51c081bf",
  1446 => x"dcc47ec1",
  1447 => x"87e1e287",
  1448 => x"58a6e4c0",
  1449 => x"c087dae2",
  1450 => x"c058a6e8",
  1451 => x"c005a8ec",
  1452 => x"e4c087cb",
  1453 => x"e0c048a6",
  1454 => x"c4c07866",
  1455 => x"cddfff87",
  1456 => x"4966c487",
  1457 => x"c0c191cb",
  1458 => x"80714866",
  1459 => x"4a6e7e70",
  1460 => x"496e82c8",
  1461 => x"e0c081ca",
  1462 => x"e4c05166",
  1463 => x"81c14966",
  1464 => x"8966e0c0",
  1465 => x"307148c1",
  1466 => x"89c14970",
  1467 => x"c37a9771",
  1468 => x"49bfedca",
  1469 => x"2966e0c0",
  1470 => x"484a6a97",
  1471 => x"f0c09871",
  1472 => x"496e58a6",
  1473 => x"4d6981c4",
  1474 => x"d84866dc",
  1475 => x"c002a866",
  1476 => x"a6d887c8",
  1477 => x"c078c048",
  1478 => x"a6d887c5",
  1479 => x"d878c148",
  1480 => x"e0c01e66",
  1481 => x"ff49751e",
  1482 => x"c887e7de",
  1483 => x"c04c7086",
  1484 => x"c106acb7",
  1485 => x"857487d4",
  1486 => x"7449e0c0",
  1487 => x"c14b7589",
  1488 => x"714ac4e1",
  1489 => x"87e0e5fe",
  1490 => x"e8c085c2",
  1491 => x"80c14866",
  1492 => x"58a6ecc0",
  1493 => x"4966ecc0",
  1494 => x"a97081c1",
  1495 => x"87c8c002",
  1496 => x"c048a6d8",
  1497 => x"87c5c078",
  1498 => x"c148a6d8",
  1499 => x"1e66d878",
  1500 => x"c049a4c2",
  1501 => x"887148e0",
  1502 => x"751e4970",
  1503 => x"d1ddff49",
  1504 => x"c086c887",
  1505 => x"ff01a8b7",
  1506 => x"e8c087c0",
  1507 => x"d1c00266",
  1508 => x"c9496e87",
  1509 => x"66e8c081",
  1510 => x"c1486e51",
  1511 => x"c078e6cc",
  1512 => x"496e87cc",
  1513 => x"51c281c9",
  1514 => x"efc2486e",
  1515 => x"7ec178e8",
  1516 => x"ff87c6c0",
  1517 => x"7087c7dc",
  1518 => x"c0026e4c",
  1519 => x"66c487f5",
  1520 => x"a866c848",
  1521 => x"87cbc004",
  1522 => x"c14866c4",
  1523 => x"58a6c880",
  1524 => x"c887e0c0",
  1525 => x"88c14866",
  1526 => x"c058a6cc",
  1527 => x"c6c187d5",
  1528 => x"c8c005ac",
  1529 => x"4866cc87",
  1530 => x"a6d080c1",
  1531 => x"cddbff58",
  1532 => x"d04c7087",
  1533 => x"80c14866",
  1534 => x"7458a6d4",
  1535 => x"cbc0029c",
  1536 => x"4866c487",
  1537 => x"a866c8c1",
  1538 => x"87fff204",
  1539 => x"87e5daff",
  1540 => x"c74866c4",
  1541 => x"e5c003a8",
  1542 => x"c0c7c387",
  1543 => x"c478c048",
  1544 => x"91cb4966",
  1545 => x"8166c0c1",
  1546 => x"6a4aa1c4",
  1547 => x"7952c04a",
  1548 => x"c14866c4",
  1549 => x"58a6c880",
  1550 => x"ff04a8c7",
  1551 => x"d0ff87db",
  1552 => x"87cce18e",
  1553 => x"1e00203a",
  1554 => x"4b711e73",
  1555 => x"87c6029b",
  1556 => x"48fcc6c3",
  1557 => x"1ec778c0",
  1558 => x"bffcc6c3",
  1559 => x"e4c11e49",
  1560 => x"c6c31edc",
  1561 => x"ee49bff8",
  1562 => x"86cc87f4",
  1563 => x"bff8c6c3",
  1564 => x"87caea49",
  1565 => x"c8029b73",
  1566 => x"dce4c187",
  1567 => x"f2e5c049",
  1568 => x"87d0e087",
  1569 => x"87d6c71e",
  1570 => x"fafe49c1",
  1571 => x"cfeafe87",
  1572 => x"02987087",
  1573 => x"f3fe87cd",
  1574 => x"987087cc",
  1575 => x"c187c402",
  1576 => x"c087c24a",
  1577 => x"059a724a",
  1578 => x"1ec087ce",
  1579 => x"49d5e3c1",
  1580 => x"87c4f1c0",
  1581 => x"87fe86c4",
  1582 => x"e3c11ec0",
  1583 => x"f0c049e0",
  1584 => x"1ec087f6",
  1585 => x"87e7d1c1",
  1586 => x"f0c04970",
  1587 => x"ccc387ea",
  1588 => x"268ef887",
  1589 => x"2044534f",
  1590 => x"6c696166",
  1591 => x"002e6465",
  1592 => x"746f6f42",
  1593 => x"2e676e69",
  1594 => x"1e002e2e",
  1595 => x"87d2e8c0",
  1596 => x"87faf3c0",
  1597 => x"4f2687f6",
  1598 => x"fcc6c31e",
  1599 => x"c378c048",
  1600 => x"c048f8c6",
  1601 => x"87fcfd78",
  1602 => x"48c087e1",
  1603 => x"20804f26",
  1604 => x"74697845",
  1605 => x"42208000",
  1606 => x"006b6361",
  1607 => x"000012d6",
  1608 => x"000031d1",
  1609 => x"d6000000",
  1610 => x"ef000012",
  1611 => x"00000031",
  1612 => x"12d60000",
  1613 => x"320d0000",
  1614 => x"00000000",
  1615 => x"0012d600",
  1616 => x"00322b00",
  1617 => x"00000000",
  1618 => x"000012d6",
  1619 => x"00003249",
  1620 => x"d6000000",
  1621 => x"67000012",
  1622 => x"00000032",
  1623 => x"12d60000",
  1624 => x"32850000",
  1625 => x"00000000",
  1626 => x"0012d600",
  1627 => x"00000000",
  1628 => x"00000000",
  1629 => x"0000135a",
  1630 => x"00000000",
  1631 => x"4c000000",
  1632 => x"2064616f",
  1633 => x"1e002e2a",
  1634 => x"c048f0fe",
  1635 => x"7909cd78",
  1636 => x"1e4f2609",
  1637 => x"bff0fe1e",
  1638 => x"2626487e",
  1639 => x"f0fe1e4f",
  1640 => x"2678c148",
  1641 => x"f0fe1e4f",
  1642 => x"2678c048",
  1643 => x"4a711e4f",
  1644 => x"265252c0",
  1645 => x"5b5e0e4f",
  1646 => x"f40e5d5c",
  1647 => x"974d7186",
  1648 => x"a5c17e6d",
  1649 => x"486c974c",
  1650 => x"6e58a6c8",
  1651 => x"a866c448",
  1652 => x"ff87c505",
  1653 => x"87e6c048",
  1654 => x"c287caff",
  1655 => x"6c9749a5",
  1656 => x"4ba3714b",
  1657 => x"974b6b97",
  1658 => x"486e7e6c",
  1659 => x"a6c880c1",
  1660 => x"cc98c758",
  1661 => x"977058a6",
  1662 => x"87e1fe7c",
  1663 => x"8ef44873",
  1664 => x"4c264d26",
  1665 => x"4f264b26",
  1666 => x"5c5b5e0e",
  1667 => x"7186f40e",
  1668 => x"4a66d84c",
  1669 => x"c29affc3",
  1670 => x"6c974ba4",
  1671 => x"49a17349",
  1672 => x"6c975172",
  1673 => x"c1486e7e",
  1674 => x"58a6c880",
  1675 => x"a6cc98c7",
  1676 => x"f4547058",
  1677 => x"87caff8e",
  1678 => x"e8fd1e1e",
  1679 => x"4abfe087",
  1680 => x"c0e0c049",
  1681 => x"87cb0299",
  1682 => x"cac31e72",
  1683 => x"f7fe49e3",
  1684 => x"fc86c487",
  1685 => x"7e7087fd",
  1686 => x"2687c2fd",
  1687 => x"c31e4f26",
  1688 => x"fd49e3ca",
  1689 => x"e8c187c7",
  1690 => x"dafc49f8",
  1691 => x"87d0c587",
  1692 => x"5e0e4f26",
  1693 => x"0e5d5c5b",
  1694 => x"bfc2cbc3",
  1695 => x"c6ebc14a",
  1696 => x"724c49bf",
  1697 => x"fc4d71bc",
  1698 => x"4bc087db",
  1699 => x"99d04974",
  1700 => x"7587d502",
  1701 => x"7199d049",
  1702 => x"c11ec01e",
  1703 => x"734acff1",
  1704 => x"c0491282",
  1705 => x"86c887e4",
  1706 => x"832d2cc1",
  1707 => x"ff04abc8",
  1708 => x"e8fb87da",
  1709 => x"c6ebc187",
  1710 => x"c2cbc348",
  1711 => x"4d2678bf",
  1712 => x"4b264c26",
  1713 => x"00004f26",
  1714 => x"ff1e0000",
  1715 => x"e1c848d0",
  1716 => x"48d4ff78",
  1717 => x"66c478c5",
  1718 => x"c387c302",
  1719 => x"66c878e0",
  1720 => x"ff87c602",
  1721 => x"f0c348d4",
  1722 => x"48d4ff78",
  1723 => x"d0ff7871",
  1724 => x"78e1c848",
  1725 => x"2678e0c0",
  1726 => x"5b5e0e4f",
  1727 => x"4c710e5c",
  1728 => x"49e3cac3",
  1729 => x"7087eefa",
  1730 => x"aab7c04a",
  1731 => x"87e3c204",
  1732 => x"05aae0c3",
  1733 => x"eec187c9",
  1734 => x"78c148fc",
  1735 => x"c387d4c2",
  1736 => x"c905aaf0",
  1737 => x"f8eec187",
  1738 => x"c178c148",
  1739 => x"eec187f5",
  1740 => x"c702bffc",
  1741 => x"c24b7287",
  1742 => x"87c2b3c0",
  1743 => x"9c744b72",
  1744 => x"c187d105",
  1745 => x"1ebff8ee",
  1746 => x"bffceec1",
  1747 => x"fd49721e",
  1748 => x"86c887f8",
  1749 => x"bff8eec1",
  1750 => x"87e0c002",
  1751 => x"b7c44973",
  1752 => x"f0c19129",
  1753 => x"4a7381cf",
  1754 => x"92c29acf",
  1755 => x"307248c1",
  1756 => x"baff4a70",
  1757 => x"98694872",
  1758 => x"87db7970",
  1759 => x"b7c44973",
  1760 => x"f0c19129",
  1761 => x"4a7381cf",
  1762 => x"92c29acf",
  1763 => x"307248c3",
  1764 => x"69484a70",
  1765 => x"c17970b0",
  1766 => x"c048fcee",
  1767 => x"f8eec178",
  1768 => x"c378c048",
  1769 => x"f849e3ca",
  1770 => x"4a7087cb",
  1771 => x"03aab7c0",
  1772 => x"c087ddfd",
  1773 => x"87c8fc48",
  1774 => x"00000000",
  1775 => x"00000000",
  1776 => x"724ac01e",
  1777 => x"c191c449",
  1778 => x"c081cff0",
  1779 => x"d082c179",
  1780 => x"ee04aab7",
  1781 => x"0e4f2687",
  1782 => x"5d5c5b5e",
  1783 => x"f74d710e",
  1784 => x"4a7587c3",
  1785 => x"922ab7c4",
  1786 => x"82cff0c1",
  1787 => x"9ccf4c75",
  1788 => x"496a94c2",
  1789 => x"c32b744b",
  1790 => x"7448c29b",
  1791 => x"ff4c7030",
  1792 => x"714874bc",
  1793 => x"f67a7098",
  1794 => x"487387d3",
  1795 => x"0087effa",
  1796 => x"00000000",
  1797 => x"00000000",
  1798 => x"00000000",
  1799 => x"00000000",
  1800 => x"00000000",
  1801 => x"00000000",
  1802 => x"00000000",
  1803 => x"00000000",
  1804 => x"00000000",
  1805 => x"00000000",
  1806 => x"00000000",
  1807 => x"00000000",
  1808 => x"00000000",
  1809 => x"00000000",
  1810 => x"00000000",
  1811 => x"16000000",
  1812 => x"2e25261e",
  1813 => x"1e3e3d36",
  1814 => x"c848d0ff",
  1815 => x"487178e1",
  1816 => x"7808d4ff",
  1817 => x"ff1e4f26",
  1818 => x"e1c848d0",
  1819 => x"ff487178",
  1820 => x"c47808d4",
  1821 => x"d4ff4866",
  1822 => x"4f267808",
  1823 => x"c44a711e",
  1824 => x"721e4966",
  1825 => x"87deff49",
  1826 => x"c048d0ff",
  1827 => x"262678e0",
  1828 => x"4a711e4f",
  1829 => x"c11e66c4",
  1830 => x"ff49a2e0",
  1831 => x"66c887c8",
  1832 => x"29b7c849",
  1833 => x"7148d4ff",
  1834 => x"48d0ff78",
  1835 => x"2678e0c0",
  1836 => x"711e4f26",
  1837 => x"49da1e4a",
  1838 => x"c887ebfe",
  1839 => x"c849bf66",
  1840 => x"80c44866",
  1841 => x"c858a6cc",
  1842 => x"d4ff29b7",
  1843 => x"c8787148",
  1844 => x"c849bf66",
  1845 => x"787129b7",
  1846 => x"c048d0ff",
  1847 => x"262678e0",
  1848 => x"d4ff1e4f",
  1849 => x"7affc34a",
  1850 => x"c848d0ff",
  1851 => x"7ade78e1",
  1852 => x"bfedcac3",
  1853 => x"c848497a",
  1854 => x"717a7028",
  1855 => x"7028d048",
  1856 => x"d848717a",
  1857 => x"ff7a7028",
  1858 => x"e0c048d0",
  1859 => x"0e4f2678",
  1860 => x"5d5c5b5e",
  1861 => x"c34c710e",
  1862 => x"4dbfedca",
  1863 => x"d02b744b",
  1864 => x"83c19b66",
  1865 => x"04ab66d4",
  1866 => x"4bc087c2",
  1867 => x"66d04a74",
  1868 => x"ff317249",
  1869 => x"739975b9",
  1870 => x"70307248",
  1871 => x"b071484a",
  1872 => x"58f1cac3",
  1873 => x"2687dafe",
  1874 => x"264c264d",
  1875 => x"1e4f264b",
  1876 => x"c848d0ff",
  1877 => x"487178c9",
  1878 => x"7808d4ff",
  1879 => x"711e4f26",
  1880 => x"87eb494a",
  1881 => x"c848d0ff",
  1882 => x"1e4f2678",
  1883 => x"4b711e73",
  1884 => x"bffdcac3",
  1885 => x"c287c302",
  1886 => x"d0ff87eb",
  1887 => x"78c9c848",
  1888 => x"e0c04973",
  1889 => x"48d4ffb1",
  1890 => x"cac37871",
  1891 => x"78c048f1",
  1892 => x"c50266c8",
  1893 => x"49ffc387",
  1894 => x"49c087c2",
  1895 => x"59f9cac3",
  1896 => x"c60266cc",
  1897 => x"d5d5c587",
  1898 => x"cf87c44a",
  1899 => x"c34affff",
  1900 => x"c35afdca",
  1901 => x"c148fdca",
  1902 => x"2687c478",
  1903 => x"264c264d",
  1904 => x"0e4f264b",
  1905 => x"5d5c5b5e",
  1906 => x"c34a710e",
  1907 => x"4cbff9ca",
  1908 => x"cb029a72",
  1909 => x"91c84987",
  1910 => x"4be1f5c1",
  1911 => x"87c48371",
  1912 => x"4be1f9c1",
  1913 => x"49134dc0",
  1914 => x"cac39974",
  1915 => x"ffb9bff5",
  1916 => x"787148d4",
  1917 => x"852cb7c1",
  1918 => x"04adb7c8",
  1919 => x"cac387e8",
  1920 => x"c848bff1",
  1921 => x"f5cac380",
  1922 => x"87effe58",
  1923 => x"711e731e",
  1924 => x"9a4a134b",
  1925 => x"7287cb02",
  1926 => x"87e7fe49",
  1927 => x"059a4a13",
  1928 => x"dafe87f5",
  1929 => x"cac31e87",
  1930 => x"c349bff1",
  1931 => x"c148f1ca",
  1932 => x"c0c478a1",
  1933 => x"db03a9b7",
  1934 => x"48d4ff87",
  1935 => x"bff5cac3",
  1936 => x"f1cac378",
  1937 => x"cac349bf",
  1938 => x"a1c148f1",
  1939 => x"b7c0c478",
  1940 => x"87e504a9",
  1941 => x"c848d0ff",
  1942 => x"fdcac378",
  1943 => x"2678c048",
  1944 => x"0000004f",
  1945 => x"00000000",
  1946 => x"00000000",
  1947 => x"00005f5f",
  1948 => x"03030000",
  1949 => x"00030300",
  1950 => x"7f7f1400",
  1951 => x"147f7f14",
  1952 => x"2e240000",
  1953 => x"123a6b6b",
  1954 => x"366a4c00",
  1955 => x"32566c18",
  1956 => x"4f7e3000",
  1957 => x"683a7759",
  1958 => x"04000040",
  1959 => x"00000307",
  1960 => x"1c000000",
  1961 => x"0041633e",
  1962 => x"41000000",
  1963 => x"001c3e63",
  1964 => x"3e2a0800",
  1965 => x"2a3e1c1c",
  1966 => x"08080008",
  1967 => x"08083e3e",
  1968 => x"80000000",
  1969 => x"000060e0",
  1970 => x"08080000",
  1971 => x"08080808",
  1972 => x"00000000",
  1973 => x"00006060",
  1974 => x"30604000",
  1975 => x"03060c18",
  1976 => x"7f3e0001",
  1977 => x"3e7f4d59",
  1978 => x"06040000",
  1979 => x"00007f7f",
  1980 => x"63420000",
  1981 => x"464f5971",
  1982 => x"63220000",
  1983 => x"367f4949",
  1984 => x"161c1800",
  1985 => x"107f7f13",
  1986 => x"67270000",
  1987 => x"397d4545",
  1988 => x"7e3c0000",
  1989 => x"3079494b",
  1990 => x"01010000",
  1991 => x"070f7971",
  1992 => x"7f360000",
  1993 => x"367f4949",
  1994 => x"4f060000",
  1995 => x"1e3f6949",
  1996 => x"00000000",
  1997 => x"00006666",
  1998 => x"80000000",
  1999 => x"000066e6",
  2000 => x"08080000",
  2001 => x"22221414",
  2002 => x"14140000",
  2003 => x"14141414",
  2004 => x"22220000",
  2005 => x"08081414",
  2006 => x"03020000",
  2007 => x"060f5951",
  2008 => x"417f3e00",
  2009 => x"1e1f555d",
  2010 => x"7f7e0000",
  2011 => x"7e7f0909",
  2012 => x"7f7f0000",
  2013 => x"367f4949",
  2014 => x"3e1c0000",
  2015 => x"41414163",
  2016 => x"7f7f0000",
  2017 => x"1c3e6341",
  2018 => x"7f7f0000",
  2019 => x"41414949",
  2020 => x"7f7f0000",
  2021 => x"01010909",
  2022 => x"7f3e0000",
  2023 => x"7a7b4941",
  2024 => x"7f7f0000",
  2025 => x"7f7f0808",
  2026 => x"41000000",
  2027 => x"00417f7f",
  2028 => x"60200000",
  2029 => x"3f7f4040",
  2030 => x"087f7f00",
  2031 => x"4163361c",
  2032 => x"7f7f0000",
  2033 => x"40404040",
  2034 => x"067f7f00",
  2035 => x"7f7f060c",
  2036 => x"067f7f00",
  2037 => x"7f7f180c",
  2038 => x"7f3e0000",
  2039 => x"3e7f4141",
  2040 => x"7f7f0000",
  2041 => x"060f0909",
  2042 => x"417f3e00",
  2043 => x"407e7f61",
  2044 => x"7f7f0000",
  2045 => x"667f1909",
  2046 => x"6f260000",
  2047 => x"327b594d",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
