//-------------------------------------------------------------------------------------------------
module rom
//-------------------------------------------------------------------------------------------------
#
(
	parameter addrbits = 0,
	parameter init_file = ""
)
(
	input  wire clock,
	input  wire ce,
	output reg  [7:0] q,
	input  wire [addrbits-1:0] a
);
//-------------------------------------------------------------------------------------------------

reg[7:0] rom[(2**addrbits)-1:0];
initial $readmemh(init_file, rom, 0);

always @(posedge clock) if(ce) q <= rom[a];

//-------------------------------------------------------------------------------------------------
endmodule
//-------------------------------------------------------------------------------------------------
