library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom2 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"4b264c26",
     1 => x"711e4f26",
     2 => x"d2eec24a",
     3 => x"d2eec25a",
     4 => x"4978c748",
     5 => x"2687ddfe",
     6 => x"1e731e4f",
     7 => x"b7c04a71",
     8 => x"87d303aa",
     9 => x"bff0cec2",
    10 => x"c187c405",
    11 => x"c087c24b",
    12 => x"f4cec24b",
    13 => x"c287c45b",
    14 => x"c25af4ce",
    15 => x"4abff0ce",
    16 => x"c0c19ac1",
    17 => x"e8ec49a2",
    18 => x"c248fc87",
    19 => x"78bff0ce",
    20 => x"1e87effe",
    21 => x"66c44a71",
    22 => x"e949721e",
    23 => x"262687f5",
    24 => x"cec21e4f",
    25 => x"e649bff0",
    26 => x"eec287cf",
    27 => x"bfe848c6",
    28 => x"c2eec278",
    29 => x"78bfec48",
    30 => x"bfc6eec2",
    31 => x"ffc3494a",
    32 => x"2ab7c899",
    33 => x"b0714872",
    34 => x"58ceeec2",
    35 => x"5e0e4f26",
    36 => x"0e5d5c5b",
    37 => x"c8ff4b71",
    38 => x"c1eec287",
    39 => x"7350c048",
    40 => x"87f5e549",
    41 => x"c24c4970",
    42 => x"49eecb9c",
    43 => x"7087c9cc",
    44 => x"eec24d49",
    45 => x"05bf97c1",
    46 => x"d087e2c1",
    47 => x"eec24966",
    48 => x"0599bfca",
    49 => x"66d487d6",
    50 => x"c2eec249",
    51 => x"cb0599bf",
    52 => x"e5497387",
    53 => x"987087c3",
    54 => x"87c1c102",
    55 => x"c0fe4cc1",
    56 => x"cb497587",
    57 => x"987087de",
    58 => x"c287c602",
    59 => x"c148c1ee",
    60 => x"c1eec250",
    61 => x"c005bf97",
    62 => x"eec287e3",
    63 => x"d049bfca",
    64 => x"ff059966",
    65 => x"eec287d6",
    66 => x"d449bfc2",
    67 => x"ff059966",
    68 => x"497387ca",
    69 => x"7087c2e4",
    70 => x"fffe0598",
    71 => x"fb487487",
    72 => x"5e0e87dc",
    73 => x"0e5d5c5b",
    74 => x"4dc086f4",
    75 => x"7ebfec4c",
    76 => x"c248a6c4",
    77 => x"78bfceee",
    78 => x"1ec01ec1",
    79 => x"cdfd49c7",
    80 => x"7086c887",
    81 => x"87cd0298",
    82 => x"ccfb49ff",
    83 => x"49dac187",
    84 => x"c187c6e3",
    85 => x"c1eec24d",
    86 => x"c302bf97",
    87 => x"87eed587",
    88 => x"bfc6eec2",
    89 => x"f0cec24b",
    90 => x"d9c105bf",
    91 => x"48a6c487",
    92 => x"78c0c0c8",
    93 => x"7edccec2",
    94 => x"49bf976e",
    95 => x"80c1486e",
    96 => x"e2717e70",
    97 => x"987087d3",
    98 => x"c487c302",
    99 => x"66c4b366",
   100 => x"28b7c148",
   101 => x"7058a6c8",
   102 => x"dbff0598",
   103 => x"49fdc387",
   104 => x"c387f6e1",
   105 => x"f0e149fa",
   106 => x"c3497387",
   107 => x"1e7199ff",
   108 => x"defa49c0",
   109 => x"c8497387",
   110 => x"1e7129b7",
   111 => x"d2fa49c1",
   112 => x"c586c887",
   113 => x"eec287ff",
   114 => x"9b4bbfca",
   115 => x"c287dd02",
   116 => x"49bfecce",
   117 => x"7087edc7",
   118 => x"87c40598",
   119 => x"87d24bc0",
   120 => x"c749e0c2",
   121 => x"cec287d2",
   122 => x"87c658f0",
   123 => x"48eccec2",
   124 => x"497378c0",
   125 => x"cd0599c2",
   126 => x"49ebc387",
   127 => x"7087dae0",
   128 => x"0299c249",
   129 => x"4cfb87c2",
   130 => x"99c14973",
   131 => x"c387cd05",
   132 => x"c4e049f4",
   133 => x"c2497087",
   134 => x"87c20299",
   135 => x"49734cfa",
   136 => x"ce0599c8",
   137 => x"49f5c387",
   138 => x"87eddfff",
   139 => x"99c24970",
   140 => x"c287d502",
   141 => x"02bfd2ee",
   142 => x"c14887ca",
   143 => x"d6eec288",
   144 => x"87c2c058",
   145 => x"4dc14cff",
   146 => x"99c44973",
   147 => x"c387ce05",
   148 => x"dfff49f2",
   149 => x"497087c3",
   150 => x"dc0299c2",
   151 => x"d2eec287",
   152 => x"c7487ebf",
   153 => x"c003a8b7",
   154 => x"486e87cb",
   155 => x"eec280c1",
   156 => x"c2c058d6",
   157 => x"c14cfe87",
   158 => x"49fdc34d",
   159 => x"87d9deff",
   160 => x"99c24970",
   161 => x"87d5c002",
   162 => x"bfd2eec2",
   163 => x"87c9c002",
   164 => x"48d2eec2",
   165 => x"c2c078c0",
   166 => x"c14cfd87",
   167 => x"49fac34d",
   168 => x"87f5ddff",
   169 => x"99c24970",
   170 => x"87d9c002",
   171 => x"bfd2eec2",
   172 => x"a8b7c748",
   173 => x"87c9c003",
   174 => x"48d2eec2",
   175 => x"c2c078c7",
   176 => x"c14cfc87",
   177 => x"acb7c04d",
   178 => x"87d1c003",
   179 => x"c14a66c4",
   180 => x"026a82d8",
   181 => x"6a87c6c0",
   182 => x"7349744b",
   183 => x"c31ec00f",
   184 => x"dac11ef0",
   185 => x"87e6f649",
   186 => x"987086c8",
   187 => x"87e2c002",
   188 => x"c248a6c8",
   189 => x"78bfd2ee",
   190 => x"cb4966c8",
   191 => x"4866c491",
   192 => x"7e708071",
   193 => x"c002bf6e",
   194 => x"bf6e87c8",
   195 => x"4966c84b",
   196 => x"9d750f73",
   197 => x"87c8c002",
   198 => x"bfd2eec2",
   199 => x"87d4f249",
   200 => x"bff4cec2",
   201 => x"87ddc002",
   202 => x"87d8c249",
   203 => x"c0029870",
   204 => x"eec287d3",
   205 => x"f149bfd2",
   206 => x"49c087fa",
   207 => x"c287daf3",
   208 => x"c048f4ce",
   209 => x"f28ef478",
   210 => x"5e0e87f4",
   211 => x"0e5d5c5b",
   212 => x"c24c711e",
   213 => x"49bfceee",
   214 => x"4da1cdc1",
   215 => x"6981d1c1",
   216 => x"029c747e",
   217 => x"a5c487cf",
   218 => x"c27b744b",
   219 => x"49bfceee",
   220 => x"6e87d3f2",
   221 => x"059c747b",
   222 => x"4bc087c4",
   223 => x"4bc187c2",
   224 => x"d4f24973",
   225 => x"0266d487",
   226 => x"c04987c8",
   227 => x"4a7087ea",
   228 => x"4ac087c2",
   229 => x"5af8cec2",
   230 => x"87e2f126",
   231 => x"14111258",
   232 => x"231c1b1d",
   233 => x"9491595a",
   234 => x"f4ebf2f5",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"ff4a711e",
   239 => x"7249bfc8",
   240 => x"4f2648a1",
   241 => x"bfc8ff1e",
   242 => x"c0c0fe89",
   243 => x"a9c0c0c0",
   244 => x"c087c401",
   245 => x"c187c24a",
   246 => x"2648724a",
   247 => x"5b5e0e4f",
   248 => x"710e5d5c",
   249 => x"4cd4ff4b",
   250 => x"c04866d0",
   251 => x"ff49d678",
   252 => x"c387e6da",
   253 => x"496c7cff",
   254 => x"7199ffc3",
   255 => x"f0c3494d",
   256 => x"a9e0c199",
   257 => x"c387cb05",
   258 => x"486c7cff",
   259 => x"66d098c3",
   260 => x"ffc37808",
   261 => x"494a6c7c",
   262 => x"ffc331c8",
   263 => x"714a6c7c",
   264 => x"c84972b2",
   265 => x"7cffc331",
   266 => x"b2714a6c",
   267 => x"31c84972",
   268 => x"6c7cffc3",
   269 => x"ffb2714a",
   270 => x"e0c048d0",
   271 => x"029b7378",
   272 => x"7b7287c2",
   273 => x"4d264875",
   274 => x"4b264c26",
   275 => x"261e4f26",
   276 => x"5b5e0e4f",
   277 => x"86f80e5c",
   278 => x"a6c81e76",
   279 => x"87fdfd49",
   280 => x"4b7086c4",
   281 => x"a8c2486e",
   282 => x"87f0c203",
   283 => x"f0c34a73",
   284 => x"aad0c19a",
   285 => x"c187c702",
   286 => x"c205aae0",
   287 => x"497387de",
   288 => x"c30299c8",
   289 => x"87c6ff87",
   290 => x"9cc34c73",
   291 => x"c105acc2",
   292 => x"66c487c2",
   293 => x"7131c949",
   294 => x"4a66c41e",
   295 => x"eec292d4",
   296 => x"817249d6",
   297 => x"87c7d4fe",
   298 => x"d7ff49d8",
   299 => x"c0c887eb",
   300 => x"c6ddc21e",
   301 => x"e2f0fd49",
   302 => x"48d0ff87",
   303 => x"c278e0c0",
   304 => x"cc1ec6dd",
   305 => x"92d44a66",
   306 => x"49d6eec2",
   307 => x"d2fe8172",
   308 => x"86cc87da",
   309 => x"c105acc1",
   310 => x"66c487c2",
   311 => x"7131c949",
   312 => x"4a66c41e",
   313 => x"eec292d4",
   314 => x"817249d6",
   315 => x"87ffd2fe",
   316 => x"1ec6ddc2",
   317 => x"d44a66c8",
   318 => x"d6eec292",
   319 => x"fe817249",
   320 => x"d787e6d0",
   321 => x"d0d6ff49",
   322 => x"1ec0c887",
   323 => x"49c6ddc2",
   324 => x"87f1eefd",
   325 => x"d0ff86cc",
   326 => x"78e0c048",
   327 => x"e7fc8ef8",
   328 => x"5b5e0e87",
   329 => x"1e0e5d5c",
   330 => x"d4ff4d71",
   331 => x"7e66d44c",
   332 => x"a8b7c348",
   333 => x"c087c506",
   334 => x"87e2c148",
   335 => x"e0fe4975",
   336 => x"1e7587fe",
   337 => x"d44b66c4",
   338 => x"d6eec293",
   339 => x"fe497383",
   340 => x"c887facb",
   341 => x"ff4b6b83",
   342 => x"e1c848d0",
   343 => x"737cdd78",
   344 => x"99ffc349",
   345 => x"49737c71",
   346 => x"c329b7c8",
   347 => x"7c7199ff",
   348 => x"b7d04973",
   349 => x"99ffc329",
   350 => x"49737c71",
   351 => x"7129b7d8",
   352 => x"7c7cc07c",
   353 => x"7c7c7c7c",
   354 => x"7c7c7c7c",
   355 => x"e0c07c7c",
   356 => x"1e66c478",
   357 => x"d4ff49dc",
   358 => x"86c887e4",
   359 => x"fa264873",
   360 => x"5e0e87e4",
   361 => x"0e5d5c5b",
   362 => x"ff7e711e",
   363 => x"1e6e4bd4",
   364 => x"49feeec2",
   365 => x"87d5cafe",
   366 => x"4d7086c4",
   367 => x"c3c3029d",
   368 => x"c6efc287",
   369 => x"496e4cbf",
   370 => x"87f4defe",
   371 => x"c848d0ff",
   372 => x"d6c178c5",
   373 => x"154ac07b",
   374 => x"c082c17b",
   375 => x"04aab7e0",
   376 => x"d0ff87f5",
   377 => x"c878c448",
   378 => x"d3c178c5",
   379 => x"c47bc17b",
   380 => x"029c7478",
   381 => x"c287fcc1",
   382 => x"c87ec6dd",
   383 => x"c08c4dc0",
   384 => x"c603acb7",
   385 => x"a4c0c887",
   386 => x"c24cc04d",
   387 => x"bf97f7e9",
   388 => x"0299d049",
   389 => x"1ec087d2",
   390 => x"49feeec2",
   391 => x"87c9ccfe",
   392 => x"497086c4",
   393 => x"87efc04a",
   394 => x"1ec6ddc2",
   395 => x"49feeec2",
   396 => x"87f5cbfe",
   397 => x"497086c4",
   398 => x"48d0ff4a",
   399 => x"c178c5c8",
   400 => x"976e7bd4",
   401 => x"486e7bbf",
   402 => x"7e7080c1",
   403 => x"ff058dc1",
   404 => x"d0ff87f0",
   405 => x"7278c448",
   406 => x"87c5059a",
   407 => x"e5c048c0",
   408 => x"c21ec187",
   409 => x"fe49feee",
   410 => x"c487ddc9",
   411 => x"059c7486",
   412 => x"ff87c4fe",
   413 => x"c5c848d0",
   414 => x"7bd3c178",
   415 => x"78c47bc0",
   416 => x"87c248c1",
   417 => x"262648c0",
   418 => x"264c264d",
   419 => x"0e4f264b",
   420 => x"0e5c5b5e",
   421 => x"66cc4b71",
   422 => x"4c87d802",
   423 => x"028cf0c0",
   424 => x"4a7487d8",
   425 => x"d1028ac1",
   426 => x"cd028a87",
   427 => x"c9028a87",
   428 => x"7387d787",
   429 => x"87eafb49",
   430 => x"1e7487d0",
   431 => x"e0f949c0",
   432 => x"731e7487",
   433 => x"87d9f949",
   434 => x"fcfe86c8",
   435 => x"c21e0087",
   436 => x"49bfdcdc",
   437 => x"dcc2b9c1",
   438 => x"d4ff59e0",
   439 => x"78ffc348",
   440 => x"c848d0ff",
   441 => x"d4ff78e1",
   442 => x"c478c148",
   443 => x"ff787131",
   444 => x"e0c048d0",
   445 => x"1e4f2678",
   446 => x"1ed0dcc2",
   447 => x"49feeec2",
   448 => x"87c9c5fe",
   449 => x"987086c4",
   450 => x"ff87c302",
   451 => x"4f2687c0",
   452 => x"484b3531",
   453 => x"2020205a",
   454 => x"00474643",
   455 => x"00000000",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
