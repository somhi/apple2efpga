
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom1 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"f4",x"d3",x"c3",x"87"),
    12 => (x"86",x"c0",x"c6",x"4e"),
    13 => (x"49",x"f4",x"d3",x"c3"),
    14 => (x"48",x"e0",x"f9",x"c2"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"ed",x"e2"),
    19 => (x"1e",x"87",x"fc",x"98"),
    20 => (x"1e",x"73",x"1e",x"72"),
    21 => (x"02",x"11",x"48",x"12"),
    22 => (x"c3",x"4b",x"87",x"ca"),
    23 => (x"73",x"9b",x"98",x"df"),
    24 => (x"87",x"f0",x"02",x"88"),
    25 => (x"4a",x"26",x"4b",x"26"),
    26 => (x"73",x"1e",x"4f",x"26"),
    27 => (x"c1",x"1e",x"72",x"1e"),
    28 => (x"87",x"ca",x"04",x"8b"),
    29 => (x"02",x"11",x"48",x"12"),
    30 => (x"02",x"88",x"87",x"c4"),
    31 => (x"4a",x"26",x"87",x"f1"),
    32 => (x"4f",x"26",x"4b",x"26"),
    33 => (x"73",x"1e",x"74",x"1e"),
    34 => (x"c1",x"1e",x"72",x"1e"),
    35 => (x"87",x"d0",x"04",x"8b"),
    36 => (x"02",x"11",x"48",x"12"),
    37 => (x"c3",x"4c",x"87",x"ca"),
    38 => (x"74",x"9c",x"98",x"df"),
    39 => (x"87",x"eb",x"02",x"88"),
    40 => (x"4b",x"26",x"4a",x"26"),
    41 => (x"4f",x"26",x"4c",x"26"),
    42 => (x"81",x"48",x"73",x"1e"),
    43 => (x"c5",x"02",x"a9",x"73"),
    44 => (x"05",x"53",x"12",x"87"),
    45 => (x"4f",x"26",x"87",x"f6"),
    46 => (x"4a",x"66",x"c4",x"1e"),
    47 => (x"51",x"12",x"48",x"71"),
    48 => (x"26",x"87",x"fb",x"05"),
    49 => (x"1e",x"73",x"1e",x"4f"),
    50 => (x"c0",x"02",x"9a",x"72"),
    51 => (x"48",x"c0",x"87",x"e7"),
    52 => (x"a9",x"72",x"4b",x"c1"),
    53 => (x"72",x"87",x"d1",x"06"),
    54 => (x"87",x"c9",x"06",x"82"),
    55 => (x"a9",x"72",x"83",x"73"),
    56 => (x"c3",x"87",x"f4",x"01"),
    57 => (x"3a",x"b2",x"c1",x"87"),
    58 => (x"89",x"03",x"a9",x"72"),
    59 => (x"c1",x"07",x"80",x"73"),
    60 => (x"f3",x"05",x"2b",x"2a"),
    61 => (x"26",x"4b",x"26",x"87"),
    62 => (x"1e",x"75",x"1e",x"4f"),
    63 => (x"b7",x"71",x"4d",x"c4"),
    64 => (x"b9",x"ff",x"04",x"a1"),
    65 => (x"bd",x"c3",x"81",x"c1"),
    66 => (x"a2",x"b7",x"72",x"07"),
    67 => (x"c1",x"ba",x"ff",x"04"),
    68 => (x"07",x"bd",x"c1",x"82"),
    69 => (x"c1",x"87",x"ee",x"fe"),
    70 => (x"b8",x"ff",x"04",x"2d"),
    71 => (x"2d",x"07",x"80",x"c1"),
    72 => (x"c1",x"b9",x"ff",x"04"),
    73 => (x"4d",x"26",x"07",x"81"),
    74 => (x"11",x"1e",x"4f",x"26"),
    75 => (x"08",x"d4",x"ff",x"48"),
    76 => (x"48",x"66",x"c4",x"78"),
    77 => (x"a6",x"c8",x"88",x"c1"),
    78 => (x"05",x"98",x"70",x"58"),
    79 => (x"4f",x"26",x"87",x"ed"),
    80 => (x"48",x"d4",x"ff",x"1e"),
    81 => (x"68",x"78",x"ff",x"c3"),
    82 => (x"48",x"66",x"c4",x"51"),
    83 => (x"a6",x"c8",x"88",x"c1"),
    84 => (x"05",x"98",x"70",x"58"),
    85 => (x"4f",x"26",x"87",x"eb"),
    86 => (x"ff",x"1e",x"73",x"1e"),
    87 => (x"ff",x"c3",x"4b",x"d4"),
    88 => (x"c3",x"4a",x"6b",x"7b"),
    89 => (x"49",x"6b",x"7b",x"ff"),
    90 => (x"b1",x"72",x"32",x"c8"),
    91 => (x"6b",x"7b",x"ff",x"c3"),
    92 => (x"71",x"31",x"c8",x"4a"),
    93 => (x"7b",x"ff",x"c3",x"b2"),
    94 => (x"32",x"c8",x"49",x"6b"),
    95 => (x"48",x"71",x"b1",x"72"),
    96 => (x"4d",x"26",x"87",x"c4"),
    97 => (x"4b",x"26",x"4c",x"26"),
    98 => (x"5e",x"0e",x"4f",x"26"),
    99 => (x"0e",x"5d",x"5c",x"5b"),
   100 => (x"d4",x"ff",x"4a",x"71"),
   101 => (x"c3",x"49",x"72",x"4c"),
   102 => (x"7c",x"71",x"99",x"ff"),
   103 => (x"bf",x"e0",x"f9",x"c2"),
   104 => (x"d0",x"87",x"c8",x"05"),
   105 => (x"30",x"c9",x"48",x"66"),
   106 => (x"d0",x"58",x"a6",x"d4"),
   107 => (x"29",x"d8",x"49",x"66"),
   108 => (x"71",x"99",x"ff",x"c3"),
   109 => (x"49",x"66",x"d0",x"7c"),
   110 => (x"ff",x"c3",x"29",x"d0"),
   111 => (x"d0",x"7c",x"71",x"99"),
   112 => (x"29",x"c8",x"49",x"66"),
   113 => (x"71",x"99",x"ff",x"c3"),
   114 => (x"49",x"66",x"d0",x"7c"),
   115 => (x"71",x"99",x"ff",x"c3"),
   116 => (x"d0",x"49",x"72",x"7c"),
   117 => (x"99",x"ff",x"c3",x"29"),
   118 => (x"4b",x"6c",x"7c",x"71"),
   119 => (x"4d",x"ff",x"f0",x"c9"),
   120 => (x"05",x"ab",x"ff",x"c3"),
   121 => (x"ff",x"c3",x"87",x"d0"),
   122 => (x"c1",x"4b",x"6c",x"7c"),
   123 => (x"87",x"c6",x"02",x"8d"),
   124 => (x"02",x"ab",x"ff",x"c3"),
   125 => (x"48",x"73",x"87",x"f0"),
   126 => (x"1e",x"87",x"c7",x"fe"),
   127 => (x"d4",x"ff",x"49",x"c0"),
   128 => (x"78",x"ff",x"c3",x"48"),
   129 => (x"c8",x"c3",x"81",x"c1"),
   130 => (x"f1",x"04",x"a9",x"b7"),
   131 => (x"1e",x"4f",x"26",x"87"),
   132 => (x"87",x"e7",x"1e",x"73"),
   133 => (x"4b",x"df",x"f8",x"c4"),
   134 => (x"ff",x"c0",x"1e",x"c0"),
   135 => (x"49",x"f7",x"c1",x"f0"),
   136 => (x"c4",x"87",x"e7",x"fd"),
   137 => (x"05",x"a8",x"c1",x"86"),
   138 => (x"ff",x"87",x"ea",x"c0"),
   139 => (x"ff",x"c3",x"48",x"d4"),
   140 => (x"c0",x"c0",x"c1",x"78"),
   141 => (x"1e",x"c0",x"c0",x"c0"),
   142 => (x"c1",x"f0",x"e1",x"c0"),
   143 => (x"c9",x"fd",x"49",x"e9"),
   144 => (x"70",x"86",x"c4",x"87"),
   145 => (x"87",x"ca",x"05",x"98"),
   146 => (x"c3",x"48",x"d4",x"ff"),
   147 => (x"48",x"c1",x"78",x"ff"),
   148 => (x"e6",x"fe",x"87",x"cb"),
   149 => (x"05",x"8b",x"c1",x"87"),
   150 => (x"c0",x"87",x"fd",x"fe"),
   151 => (x"87",x"e6",x"fc",x"48"),
   152 => (x"ff",x"1e",x"73",x"1e"),
   153 => (x"ff",x"c3",x"48",x"d4"),
   154 => (x"c0",x"4b",x"d3",x"78"),
   155 => (x"f0",x"ff",x"c0",x"1e"),
   156 => (x"fc",x"49",x"c1",x"c1"),
   157 => (x"86",x"c4",x"87",x"d4"),
   158 => (x"ca",x"05",x"98",x"70"),
   159 => (x"48",x"d4",x"ff",x"87"),
   160 => (x"c1",x"78",x"ff",x"c3"),
   161 => (x"fd",x"87",x"cb",x"48"),
   162 => (x"8b",x"c1",x"87",x"f1"),
   163 => (x"87",x"db",x"ff",x"05"),
   164 => (x"f1",x"fb",x"48",x"c0"),
   165 => (x"5b",x"5e",x"0e",x"87"),
   166 => (x"d4",x"ff",x"0e",x"5c"),
   167 => (x"87",x"db",x"fd",x"4c"),
   168 => (x"c0",x"1e",x"ea",x"c6"),
   169 => (x"c8",x"c1",x"f0",x"e1"),
   170 => (x"87",x"de",x"fb",x"49"),
   171 => (x"a8",x"c1",x"86",x"c4"),
   172 => (x"fe",x"87",x"c8",x"02"),
   173 => (x"48",x"c0",x"87",x"ea"),
   174 => (x"fa",x"87",x"e2",x"c1"),
   175 => (x"49",x"70",x"87",x"da"),
   176 => (x"99",x"ff",x"ff",x"cf"),
   177 => (x"02",x"a9",x"ea",x"c6"),
   178 => (x"d3",x"fe",x"87",x"c8"),
   179 => (x"c1",x"48",x"c0",x"87"),
   180 => (x"ff",x"c3",x"87",x"cb"),
   181 => (x"4b",x"f1",x"c0",x"7c"),
   182 => (x"70",x"87",x"f4",x"fc"),
   183 => (x"eb",x"c0",x"02",x"98"),
   184 => (x"c0",x"1e",x"c0",x"87"),
   185 => (x"fa",x"c1",x"f0",x"ff"),
   186 => (x"87",x"de",x"fa",x"49"),
   187 => (x"98",x"70",x"86",x"c4"),
   188 => (x"c3",x"87",x"d9",x"05"),
   189 => (x"49",x"6c",x"7c",x"ff"),
   190 => (x"7c",x"7c",x"ff",x"c3"),
   191 => (x"c0",x"c1",x"7c",x"7c"),
   192 => (x"87",x"c4",x"02",x"99"),
   193 => (x"87",x"d5",x"48",x"c1"),
   194 => (x"87",x"d1",x"48",x"c0"),
   195 => (x"c4",x"05",x"ab",x"c2"),
   196 => (x"c8",x"48",x"c0",x"87"),
   197 => (x"05",x"8b",x"c1",x"87"),
   198 => (x"c0",x"87",x"fd",x"fe"),
   199 => (x"87",x"e4",x"f9",x"48"),
   200 => (x"c2",x"1e",x"73",x"1e"),
   201 => (x"c1",x"48",x"e0",x"f9"),
   202 => (x"ff",x"4b",x"c7",x"78"),
   203 => (x"78",x"c2",x"48",x"d0"),
   204 => (x"ff",x"87",x"c8",x"fb"),
   205 => (x"78",x"c3",x"48",x"d0"),
   206 => (x"e5",x"c0",x"1e",x"c0"),
   207 => (x"49",x"c0",x"c1",x"d0"),
   208 => (x"c4",x"87",x"c7",x"f9"),
   209 => (x"05",x"a8",x"c1",x"86"),
   210 => (x"c2",x"4b",x"87",x"c1"),
   211 => (x"87",x"c5",x"05",x"ab"),
   212 => (x"f9",x"c0",x"48",x"c0"),
   213 => (x"05",x"8b",x"c1",x"87"),
   214 => (x"fc",x"87",x"d0",x"ff"),
   215 => (x"f9",x"c2",x"87",x"f7"),
   216 => (x"98",x"70",x"58",x"e4"),
   217 => (x"c1",x"87",x"cd",x"05"),
   218 => (x"f0",x"ff",x"c0",x"1e"),
   219 => (x"f8",x"49",x"d0",x"c1"),
   220 => (x"86",x"c4",x"87",x"d8"),
   221 => (x"c3",x"48",x"d4",x"ff"),
   222 => (x"e0",x"c4",x"78",x"ff"),
   223 => (x"e8",x"f9",x"c2",x"87"),
   224 => (x"48",x"d0",x"ff",x"58"),
   225 => (x"d4",x"ff",x"78",x"c2"),
   226 => (x"78",x"ff",x"c3",x"48"),
   227 => (x"f5",x"f7",x"48",x"c1"),
   228 => (x"5b",x"5e",x"0e",x"87"),
   229 => (x"71",x"0e",x"5d",x"5c"),
   230 => (x"4d",x"ff",x"c3",x"4a"),
   231 => (x"75",x"4c",x"d4",x"ff"),
   232 => (x"48",x"d0",x"ff",x"7c"),
   233 => (x"75",x"78",x"c3",x"c4"),
   234 => (x"c0",x"1e",x"72",x"7c"),
   235 => (x"d8",x"c1",x"f0",x"ff"),
   236 => (x"87",x"d6",x"f7",x"49"),
   237 => (x"98",x"70",x"86",x"c4"),
   238 => (x"c0",x"87",x"c5",x"02"),
   239 => (x"87",x"f0",x"c0",x"48"),
   240 => (x"fe",x"c3",x"7c",x"75"),
   241 => (x"1e",x"c0",x"c8",x"7c"),
   242 => (x"f5",x"49",x"66",x"d4"),
   243 => (x"86",x"c4",x"87",x"dc"),
   244 => (x"7c",x"75",x"7c",x"75"),
   245 => (x"da",x"d8",x"7c",x"75"),
   246 => (x"7c",x"75",x"4b",x"e0"),
   247 => (x"05",x"99",x"49",x"6c"),
   248 => (x"8b",x"c1",x"87",x"c5"),
   249 => (x"75",x"87",x"f3",x"05"),
   250 => (x"48",x"d0",x"ff",x"7c"),
   251 => (x"48",x"c1",x"78",x"c2"),
   252 => (x"1e",x"87",x"cf",x"f6"),
   253 => (x"ff",x"4a",x"d4",x"ff"),
   254 => (x"d1",x"c4",x"48",x"d0"),
   255 => (x"7a",x"ff",x"c3",x"78"),
   256 => (x"f8",x"05",x"89",x"c1"),
   257 => (x"1e",x"4f",x"26",x"87"),
   258 => (x"4b",x"71",x"1e",x"73"),
   259 => (x"df",x"cd",x"ee",x"c5"),
   260 => (x"48",x"d4",x"ff",x"4a"),
   261 => (x"68",x"78",x"ff",x"c3"),
   262 => (x"a8",x"fe",x"c3",x"48"),
   263 => (x"c1",x"87",x"c5",x"02"),
   264 => (x"87",x"ed",x"05",x"8a"),
   265 => (x"c5",x"05",x"9a",x"72"),
   266 => (x"c0",x"48",x"c0",x"87"),
   267 => (x"9b",x"73",x"87",x"ea"),
   268 => (x"c8",x"87",x"cc",x"02"),
   269 => (x"49",x"73",x"1e",x"66"),
   270 => (x"c4",x"87",x"c5",x"f4"),
   271 => (x"c8",x"87",x"c6",x"86"),
   272 => (x"ee",x"fe",x"49",x"66"),
   273 => (x"48",x"d4",x"ff",x"87"),
   274 => (x"78",x"78",x"ff",x"c3"),
   275 => (x"c5",x"05",x"9b",x"73"),
   276 => (x"48",x"d0",x"ff",x"87"),
   277 => (x"48",x"c1",x"78",x"d0"),
   278 => (x"1e",x"87",x"eb",x"f4"),
   279 => (x"4a",x"71",x"1e",x"73"),
   280 => (x"d4",x"ff",x"4b",x"c0"),
   281 => (x"78",x"ff",x"c3",x"48"),
   282 => (x"c4",x"48",x"d0",x"ff"),
   283 => (x"d4",x"ff",x"78",x"c3"),
   284 => (x"78",x"ff",x"c3",x"48"),
   285 => (x"ff",x"c0",x"1e",x"72"),
   286 => (x"49",x"d1",x"c1",x"f0"),
   287 => (x"c4",x"87",x"cb",x"f4"),
   288 => (x"05",x"98",x"70",x"86"),
   289 => (x"c0",x"c8",x"87",x"cd"),
   290 => (x"49",x"66",x"cc",x"1e"),
   291 => (x"c4",x"87",x"f8",x"fd"),
   292 => (x"ff",x"4b",x"70",x"86"),
   293 => (x"78",x"c2",x"48",x"d0"),
   294 => (x"e9",x"f3",x"48",x"73"),
   295 => (x"5b",x"5e",x"0e",x"87"),
   296 => (x"c0",x"0e",x"5d",x"5c"),
   297 => (x"f0",x"ff",x"c0",x"1e"),
   298 => (x"f3",x"49",x"c9",x"c1"),
   299 => (x"1e",x"d2",x"87",x"dc"),
   300 => (x"49",x"e8",x"f9",x"c2"),
   301 => (x"c8",x"87",x"d0",x"fd"),
   302 => (x"c1",x"4c",x"c0",x"86"),
   303 => (x"ac",x"b7",x"d2",x"84"),
   304 => (x"c2",x"87",x"f8",x"04"),
   305 => (x"bf",x"97",x"e8",x"f9"),
   306 => (x"99",x"c0",x"c3",x"49"),
   307 => (x"05",x"a9",x"c0",x"c1"),
   308 => (x"c2",x"87",x"e7",x"c0"),
   309 => (x"bf",x"97",x"ef",x"f9"),
   310 => (x"c2",x"31",x"d0",x"49"),
   311 => (x"bf",x"97",x"f0",x"f9"),
   312 => (x"72",x"32",x"c8",x"4a"),
   313 => (x"f1",x"f9",x"c2",x"b1"),
   314 => (x"b1",x"4a",x"bf",x"97"),
   315 => (x"ff",x"cf",x"4c",x"71"),
   316 => (x"c1",x"9c",x"ff",x"ff"),
   317 => (x"c1",x"34",x"ca",x"84"),
   318 => (x"f9",x"c2",x"87",x"e7"),
   319 => (x"49",x"bf",x"97",x"f1"),
   320 => (x"99",x"c6",x"31",x"c1"),
   321 => (x"97",x"f2",x"f9",x"c2"),
   322 => (x"b7",x"c7",x"4a",x"bf"),
   323 => (x"c2",x"b1",x"72",x"2a"),
   324 => (x"bf",x"97",x"ed",x"f9"),
   325 => (x"9d",x"cf",x"4d",x"4a"),
   326 => (x"97",x"ee",x"f9",x"c2"),
   327 => (x"9a",x"c3",x"4a",x"bf"),
   328 => (x"f9",x"c2",x"32",x"ca"),
   329 => (x"4b",x"bf",x"97",x"ef"),
   330 => (x"b2",x"73",x"33",x"c2"),
   331 => (x"97",x"f0",x"f9",x"c2"),
   332 => (x"c0",x"c3",x"4b",x"bf"),
   333 => (x"2b",x"b7",x"c6",x"9b"),
   334 => (x"81",x"c2",x"b2",x"73"),
   335 => (x"30",x"71",x"48",x"c1"),
   336 => (x"48",x"c1",x"49",x"70"),
   337 => (x"4d",x"70",x"30",x"75"),
   338 => (x"84",x"c1",x"4c",x"72"),
   339 => (x"c0",x"c8",x"94",x"71"),
   340 => (x"cc",x"06",x"ad",x"b7"),
   341 => (x"b7",x"34",x"c1",x"87"),
   342 => (x"b7",x"c0",x"c8",x"2d"),
   343 => (x"f4",x"ff",x"01",x"ad"),
   344 => (x"f0",x"48",x"74",x"87"),
   345 => (x"5e",x"0e",x"87",x"dc"),
   346 => (x"0e",x"5d",x"5c",x"5b"),
   347 => (x"c2",x"c3",x"86",x"f8"),
   348 => (x"78",x"c0",x"48",x"ce"),
   349 => (x"1e",x"c6",x"fa",x"c2"),
   350 => (x"de",x"fb",x"49",x"c0"),
   351 => (x"70",x"86",x"c4",x"87"),
   352 => (x"87",x"c5",x"05",x"98"),
   353 => (x"ce",x"c9",x"48",x"c0"),
   354 => (x"c1",x"4d",x"c0",x"87"),
   355 => (x"f8",x"f9",x"c0",x"7e"),
   356 => (x"fa",x"c2",x"49",x"bf"),
   357 => (x"c8",x"71",x"4a",x"fc"),
   358 => (x"87",x"ce",x"eb",x"4b"),
   359 => (x"c2",x"05",x"98",x"70"),
   360 => (x"c0",x"7e",x"c0",x"87"),
   361 => (x"49",x"bf",x"f4",x"f9"),
   362 => (x"4a",x"d8",x"fb",x"c2"),
   363 => (x"ea",x"4b",x"c8",x"71"),
   364 => (x"98",x"70",x"87",x"f8"),
   365 => (x"c0",x"87",x"c2",x"05"),
   366 => (x"c0",x"02",x"6e",x"7e"),
   367 => (x"c1",x"c3",x"87",x"fd"),
   368 => (x"c3",x"4d",x"bf",x"cc"),
   369 => (x"bf",x"9f",x"c4",x"c2"),
   370 => (x"d6",x"c5",x"48",x"7e"),
   371 => (x"c7",x"05",x"a8",x"ea"),
   372 => (x"cc",x"c1",x"c3",x"87"),
   373 => (x"87",x"ce",x"4d",x"bf"),
   374 => (x"e9",x"ca",x"48",x"6e"),
   375 => (x"c5",x"02",x"a8",x"d5"),
   376 => (x"c7",x"48",x"c0",x"87"),
   377 => (x"fa",x"c2",x"87",x"f1"),
   378 => (x"49",x"75",x"1e",x"c6"),
   379 => (x"c4",x"87",x"ec",x"f9"),
   380 => (x"05",x"98",x"70",x"86"),
   381 => (x"48",x"c0",x"87",x"c5"),
   382 => (x"c0",x"87",x"dc",x"c7"),
   383 => (x"49",x"bf",x"f4",x"f9"),
   384 => (x"4a",x"d8",x"fb",x"c2"),
   385 => (x"e9",x"4b",x"c8",x"71"),
   386 => (x"98",x"70",x"87",x"e0"),
   387 => (x"c3",x"87",x"c8",x"05"),
   388 => (x"c1",x"48",x"ce",x"c2"),
   389 => (x"c0",x"87",x"da",x"78"),
   390 => (x"49",x"bf",x"f8",x"f9"),
   391 => (x"4a",x"fc",x"fa",x"c2"),
   392 => (x"e9",x"4b",x"c8",x"71"),
   393 => (x"98",x"70",x"87",x"c4"),
   394 => (x"87",x"c5",x"c0",x"02"),
   395 => (x"e6",x"c6",x"48",x"c0"),
   396 => (x"c4",x"c2",x"c3",x"87"),
   397 => (x"c1",x"49",x"bf",x"97"),
   398 => (x"c0",x"05",x"a9",x"d5"),
   399 => (x"c2",x"c3",x"87",x"cd"),
   400 => (x"49",x"bf",x"97",x"c5"),
   401 => (x"02",x"a9",x"ea",x"c2"),
   402 => (x"c0",x"87",x"c5",x"c0"),
   403 => (x"87",x"c7",x"c6",x"48"),
   404 => (x"97",x"c6",x"fa",x"c2"),
   405 => (x"c3",x"48",x"7e",x"bf"),
   406 => (x"c0",x"02",x"a8",x"e9"),
   407 => (x"48",x"6e",x"87",x"ce"),
   408 => (x"02",x"a8",x"eb",x"c3"),
   409 => (x"c0",x"87",x"c5",x"c0"),
   410 => (x"87",x"eb",x"c5",x"48"),
   411 => (x"97",x"d1",x"fa",x"c2"),
   412 => (x"05",x"99",x"49",x"bf"),
   413 => (x"c2",x"87",x"cc",x"c0"),
   414 => (x"bf",x"97",x"d2",x"fa"),
   415 => (x"02",x"a9",x"c2",x"49"),
   416 => (x"c0",x"87",x"c5",x"c0"),
   417 => (x"87",x"cf",x"c5",x"48"),
   418 => (x"97",x"d3",x"fa",x"c2"),
   419 => (x"c2",x"c3",x"48",x"bf"),
   420 => (x"4c",x"70",x"58",x"ca"),
   421 => (x"c3",x"88",x"c1",x"48"),
   422 => (x"c2",x"58",x"ce",x"c2"),
   423 => (x"bf",x"97",x"d4",x"fa"),
   424 => (x"c2",x"81",x"75",x"49"),
   425 => (x"bf",x"97",x"d5",x"fa"),
   426 => (x"72",x"32",x"c8",x"4a"),
   427 => (x"c6",x"c3",x"7e",x"a1"),
   428 => (x"78",x"6e",x"48",x"db"),
   429 => (x"97",x"d6",x"fa",x"c2"),
   430 => (x"a6",x"c8",x"48",x"bf"),
   431 => (x"ce",x"c2",x"c3",x"58"),
   432 => (x"d4",x"c2",x"02",x"bf"),
   433 => (x"f4",x"f9",x"c0",x"87"),
   434 => (x"fb",x"c2",x"49",x"bf"),
   435 => (x"c8",x"71",x"4a",x"d8"),
   436 => (x"87",x"d6",x"e6",x"4b"),
   437 => (x"c0",x"02",x"98",x"70"),
   438 => (x"48",x"c0",x"87",x"c5"),
   439 => (x"c3",x"87",x"f8",x"c3"),
   440 => (x"4c",x"bf",x"c6",x"c2"),
   441 => (x"5c",x"ef",x"c6",x"c3"),
   442 => (x"97",x"eb",x"fa",x"c2"),
   443 => (x"31",x"c8",x"49",x"bf"),
   444 => (x"97",x"ea",x"fa",x"c2"),
   445 => (x"49",x"a1",x"4a",x"bf"),
   446 => (x"97",x"ec",x"fa",x"c2"),
   447 => (x"32",x"d0",x"4a",x"bf"),
   448 => (x"c2",x"49",x"a1",x"72"),
   449 => (x"bf",x"97",x"ed",x"fa"),
   450 => (x"72",x"32",x"d8",x"4a"),
   451 => (x"66",x"c4",x"49",x"a1"),
   452 => (x"db",x"c6",x"c3",x"91"),
   453 => (x"c6",x"c3",x"81",x"bf"),
   454 => (x"fa",x"c2",x"59",x"e3"),
   455 => (x"4a",x"bf",x"97",x"f3"),
   456 => (x"fa",x"c2",x"32",x"c8"),
   457 => (x"4b",x"bf",x"97",x"f2"),
   458 => (x"fa",x"c2",x"4a",x"a2"),
   459 => (x"4b",x"bf",x"97",x"f4"),
   460 => (x"a2",x"73",x"33",x"d0"),
   461 => (x"f5",x"fa",x"c2",x"4a"),
   462 => (x"cf",x"4b",x"bf",x"97"),
   463 => (x"73",x"33",x"d8",x"9b"),
   464 => (x"c6",x"c3",x"4a",x"a2"),
   465 => (x"c6",x"c3",x"5a",x"e7"),
   466 => (x"c2",x"4a",x"bf",x"e3"),
   467 => (x"c3",x"92",x"74",x"8a"),
   468 => (x"72",x"48",x"e7",x"c6"),
   469 => (x"ca",x"c1",x"78",x"a1"),
   470 => (x"d8",x"fa",x"c2",x"87"),
   471 => (x"c8",x"49",x"bf",x"97"),
   472 => (x"d7",x"fa",x"c2",x"31"),
   473 => (x"a1",x"4a",x"bf",x"97"),
   474 => (x"d6",x"c2",x"c3",x"49"),
   475 => (x"d2",x"c2",x"c3",x"59"),
   476 => (x"31",x"c5",x"49",x"bf"),
   477 => (x"c9",x"81",x"ff",x"c7"),
   478 => (x"ef",x"c6",x"c3",x"29"),
   479 => (x"dd",x"fa",x"c2",x"59"),
   480 => (x"c8",x"4a",x"bf",x"97"),
   481 => (x"dc",x"fa",x"c2",x"32"),
   482 => (x"a2",x"4b",x"bf",x"97"),
   483 => (x"92",x"66",x"c4",x"4a"),
   484 => (x"c6",x"c3",x"82",x"6e"),
   485 => (x"c6",x"c3",x"5a",x"eb"),
   486 => (x"78",x"c0",x"48",x"e3"),
   487 => (x"48",x"df",x"c6",x"c3"),
   488 => (x"c3",x"78",x"a1",x"72"),
   489 => (x"c3",x"48",x"ef",x"c6"),
   490 => (x"78",x"bf",x"e3",x"c6"),
   491 => (x"48",x"f3",x"c6",x"c3"),
   492 => (x"bf",x"e7",x"c6",x"c3"),
   493 => (x"ce",x"c2",x"c3",x"78"),
   494 => (x"c9",x"c0",x"02",x"bf"),
   495 => (x"c4",x"48",x"74",x"87"),
   496 => (x"c0",x"7e",x"70",x"30"),
   497 => (x"c6",x"c3",x"87",x"c9"),
   498 => (x"c4",x"48",x"bf",x"eb"),
   499 => (x"c3",x"7e",x"70",x"30"),
   500 => (x"6e",x"48",x"d2",x"c2"),
   501 => (x"f8",x"48",x"c1",x"78"),
   502 => (x"26",x"4d",x"26",x"8e"),
   503 => (x"26",x"4b",x"26",x"4c"),
   504 => (x"5b",x"5e",x"0e",x"4f"),
   505 => (x"71",x"0e",x"5d",x"5c"),
   506 => (x"ce",x"c2",x"c3",x"4a"),
   507 => (x"87",x"cb",x"02",x"bf"),
   508 => (x"2b",x"c7",x"4b",x"72"),
   509 => (x"ff",x"c1",x"4c",x"72"),
   510 => (x"72",x"87",x"c9",x"9c"),
   511 => (x"72",x"2b",x"c8",x"4b"),
   512 => (x"9c",x"ff",x"c3",x"4c"),
   513 => (x"bf",x"db",x"c6",x"c3"),
   514 => (x"f0",x"f9",x"c0",x"83"),
   515 => (x"d9",x"02",x"ab",x"bf"),
   516 => (x"f4",x"f9",x"c0",x"87"),
   517 => (x"c6",x"fa",x"c2",x"5b"),
   518 => (x"f0",x"49",x"73",x"1e"),
   519 => (x"86",x"c4",x"87",x"fd"),
   520 => (x"c5",x"05",x"98",x"70"),
   521 => (x"c0",x"48",x"c0",x"87"),
   522 => (x"c2",x"c3",x"87",x"e6"),
   523 => (x"d2",x"02",x"bf",x"ce"),
   524 => (x"c4",x"49",x"74",x"87"),
   525 => (x"c6",x"fa",x"c2",x"91"),
   526 => (x"cf",x"4d",x"69",x"81"),
   527 => (x"ff",x"ff",x"ff",x"ff"),
   528 => (x"74",x"87",x"cb",x"9d"),
   529 => (x"c2",x"91",x"c2",x"49"),
   530 => (x"9f",x"81",x"c6",x"fa"),
   531 => (x"48",x"75",x"4d",x"69"),
   532 => (x"0e",x"87",x"c6",x"fe"),
   533 => (x"5d",x"5c",x"5b",x"5e"),
   534 => (x"4d",x"71",x"1e",x"0e"),
   535 => (x"49",x"c1",x"1e",x"c0"),
   536 => (x"c4",x"87",x"f5",x"d0"),
   537 => (x"9c",x"4c",x"70",x"86"),
   538 => (x"87",x"c2",x"c1",x"02"),
   539 => (x"4a",x"d6",x"c2",x"c3"),
   540 => (x"df",x"ff",x"49",x"75"),
   541 => (x"98",x"70",x"87",x"d9"),
   542 => (x"87",x"f2",x"c0",x"02"),
   543 => (x"49",x"75",x"4a",x"74"),
   544 => (x"df",x"ff",x"4b",x"cb"),
   545 => (x"98",x"70",x"87",x"fe"),
   546 => (x"87",x"e2",x"c0",x"02"),
   547 => (x"9c",x"74",x"1e",x"c0"),
   548 => (x"c4",x"87",x"c7",x"02"),
   549 => (x"78",x"c0",x"48",x"a6"),
   550 => (x"a6",x"c4",x"87",x"c5"),
   551 => (x"c4",x"78",x"c1",x"48"),
   552 => (x"f3",x"cf",x"49",x"66"),
   553 => (x"70",x"86",x"c4",x"87"),
   554 => (x"fe",x"05",x"9c",x"4c"),
   555 => (x"48",x"74",x"87",x"fe"),
   556 => (x"87",x"e5",x"fc",x"26"),
   557 => (x"5c",x"5b",x"5e",x"0e"),
   558 => (x"86",x"f8",x"0e",x"5d"),
   559 => (x"05",x"9b",x"4b",x"71"),
   560 => (x"48",x"c0",x"87",x"c5"),
   561 => (x"c8",x"87",x"d4",x"c2"),
   562 => (x"7d",x"c0",x"4d",x"a3"),
   563 => (x"c7",x"02",x"66",x"d8"),
   564 => (x"97",x"66",x"d8",x"87"),
   565 => (x"87",x"c5",x"05",x"bf"),
   566 => (x"fe",x"c1",x"48",x"c0"),
   567 => (x"49",x"66",x"d8",x"87"),
   568 => (x"70",x"87",x"f0",x"fd"),
   569 => (x"c1",x"02",x"6e",x"7e"),
   570 => (x"49",x"6e",x"87",x"ef"),
   571 => (x"7d",x"69",x"81",x"dc"),
   572 => (x"81",x"da",x"49",x"6e"),
   573 => (x"9f",x"4c",x"a3",x"c4"),
   574 => (x"c2",x"c3",x"7c",x"69"),
   575 => (x"d0",x"02",x"bf",x"ce"),
   576 => (x"d4",x"49",x"6e",x"87"),
   577 => (x"49",x"69",x"9f",x"81"),
   578 => (x"ff",x"ff",x"c0",x"4a"),
   579 => (x"c2",x"32",x"d0",x"9a"),
   580 => (x"72",x"4a",x"c0",x"87"),
   581 => (x"80",x"6c",x"48",x"49"),
   582 => (x"7b",x"c0",x"7c",x"70"),
   583 => (x"6c",x"49",x"a3",x"cc"),
   584 => (x"49",x"a3",x"d0",x"79"),
   585 => (x"a6",x"c4",x"79",x"c0"),
   586 => (x"d4",x"78",x"c0",x"48"),
   587 => (x"66",x"c4",x"4a",x"a3"),
   588 => (x"72",x"91",x"c8",x"49"),
   589 => (x"41",x"c0",x"49",x"a1"),
   590 => (x"66",x"c4",x"79",x"6c"),
   591 => (x"c8",x"80",x"c1",x"48"),
   592 => (x"b7",x"d0",x"58",x"a6"),
   593 => (x"e2",x"ff",x"04",x"a8"),
   594 => (x"c9",x"4a",x"6d",x"87"),
   595 => (x"c2",x"2a",x"c7",x"2a"),
   596 => (x"72",x"49",x"a3",x"d4"),
   597 => (x"c2",x"48",x"6e",x"79"),
   598 => (x"f8",x"48",x"c0",x"87"),
   599 => (x"87",x"f9",x"f9",x"8e"),
   600 => (x"5c",x"5b",x"5e",x"0e"),
   601 => (x"4c",x"71",x"0e",x"5d"),
   602 => (x"48",x"f0",x"f9",x"c0"),
   603 => (x"9c",x"74",x"78",x"ff"),
   604 => (x"87",x"ca",x"c1",x"02"),
   605 => (x"69",x"49",x"a4",x"c8"),
   606 => (x"87",x"c2",x"c1",x"02"),
   607 => (x"6c",x"4a",x"66",x"d0"),
   608 => (x"a6",x"d4",x"82",x"49"),
   609 => (x"4d",x"66",x"d0",x"5a"),
   610 => (x"ca",x"c2",x"c3",x"b9"),
   611 => (x"ba",x"ff",x"4a",x"bf"),
   612 => (x"99",x"71",x"99",x"72"),
   613 => (x"87",x"e4",x"c0",x"02"),
   614 => (x"6b",x"4b",x"a4",x"c4"),
   615 => (x"87",x"c1",x"f9",x"49"),
   616 => (x"c2",x"c3",x"7b",x"70"),
   617 => (x"6c",x"49",x"bf",x"c6"),
   618 => (x"75",x"7c",x"71",x"81"),
   619 => (x"ca",x"c2",x"c3",x"b9"),
   620 => (x"ba",x"ff",x"4a",x"bf"),
   621 => (x"99",x"71",x"99",x"72"),
   622 => (x"87",x"dc",x"ff",x"05"),
   623 => (x"d8",x"f8",x"7c",x"75"),
   624 => (x"1e",x"73",x"1e",x"87"),
   625 => (x"02",x"9b",x"4b",x"71"),
   626 => (x"a3",x"c8",x"87",x"c7"),
   627 => (x"c5",x"05",x"69",x"49"),
   628 => (x"c0",x"48",x"c0",x"87"),
   629 => (x"c6",x"c3",x"87",x"eb"),
   630 => (x"c4",x"4a",x"bf",x"df"),
   631 => (x"49",x"69",x"49",x"a3"),
   632 => (x"c2",x"c3",x"89",x"c2"),
   633 => (x"71",x"91",x"bf",x"c6"),
   634 => (x"c2",x"c3",x"4a",x"a2"),
   635 => (x"6b",x"49",x"bf",x"ca"),
   636 => (x"4a",x"a2",x"71",x"99"),
   637 => (x"72",x"1e",x"66",x"c8"),
   638 => (x"87",x"df",x"e9",x"49"),
   639 => (x"49",x"70",x"86",x"c4"),
   640 => (x"87",x"d9",x"f7",x"48"),
   641 => (x"71",x"1e",x"73",x"1e"),
   642 => (x"c7",x"02",x"9b",x"4b"),
   643 => (x"49",x"a3",x"c8",x"87"),
   644 => (x"87",x"c5",x"05",x"69"),
   645 => (x"eb",x"c0",x"48",x"c0"),
   646 => (x"df",x"c6",x"c3",x"87"),
   647 => (x"a3",x"c4",x"4a",x"bf"),
   648 => (x"c2",x"49",x"69",x"49"),
   649 => (x"c6",x"c2",x"c3",x"89"),
   650 => (x"a2",x"71",x"91",x"bf"),
   651 => (x"ca",x"c2",x"c3",x"4a"),
   652 => (x"99",x"6b",x"49",x"bf"),
   653 => (x"c8",x"4a",x"a2",x"71"),
   654 => (x"49",x"72",x"1e",x"66"),
   655 => (x"c4",x"87",x"d2",x"e5"),
   656 => (x"48",x"49",x"70",x"86"),
   657 => (x"0e",x"87",x"d6",x"f6"),
   658 => (x"5d",x"5c",x"5b",x"5e"),
   659 => (x"71",x"86",x"f8",x"0e"),
   660 => (x"48",x"a6",x"c4",x"4b"),
   661 => (x"a3",x"c8",x"78",x"ff"),
   662 => (x"c0",x"4d",x"69",x"49"),
   663 => (x"4a",x"a3",x"d4",x"4c"),
   664 => (x"91",x"c8",x"49",x"74"),
   665 => (x"69",x"49",x"a1",x"72"),
   666 => (x"48",x"66",x"d8",x"49"),
   667 => (x"7e",x"70",x"88",x"71"),
   668 => (x"01",x"a9",x"66",x"d8"),
   669 => (x"ad",x"6e",x"87",x"ca"),
   670 => (x"c8",x"87",x"c5",x"06"),
   671 => (x"4d",x"6e",x"5c",x"a6"),
   672 => (x"b7",x"d0",x"84",x"c1"),
   673 => (x"d4",x"ff",x"04",x"ac"),
   674 => (x"48",x"66",x"c4",x"87"),
   675 => (x"c8",x"f5",x"8e",x"f8"),
   676 => (x"5b",x"5e",x"0e",x"87"),
   677 => (x"ec",x"0e",x"5d",x"5c"),
   678 => (x"59",x"a6",x"c8",x"86"),
   679 => (x"c1",x"48",x"a6",x"c8"),
   680 => (x"ff",x"ff",x"ff",x"ff"),
   681 => (x"80",x"c4",x"78",x"ff"),
   682 => (x"4d",x"c0",x"78",x"ff"),
   683 => (x"66",x"c4",x"4c",x"c0"),
   684 => (x"74",x"83",x"d4",x"4b"),
   685 => (x"73",x"91",x"c8",x"49"),
   686 => (x"4a",x"75",x"49",x"a1"),
   687 => (x"a2",x"73",x"92",x"c8"),
   688 => (x"6e",x"49",x"69",x"7e"),
   689 => (x"a6",x"d4",x"89",x"bf"),
   690 => (x"05",x"ad",x"74",x"59"),
   691 => (x"a6",x"d0",x"87",x"c6"),
   692 => (x"78",x"bf",x"6e",x"48"),
   693 => (x"c0",x"48",x"66",x"d0"),
   694 => (x"cf",x"04",x"a8",x"b7"),
   695 => (x"49",x"66",x"d0",x"87"),
   696 => (x"03",x"a9",x"66",x"c8"),
   697 => (x"a6",x"d0",x"87",x"c6"),
   698 => (x"59",x"a6",x"cc",x"5c"),
   699 => (x"b7",x"d0",x"84",x"c1"),
   700 => (x"f9",x"fe",x"04",x"ac"),
   701 => (x"d0",x"85",x"c1",x"87"),
   702 => (x"fe",x"04",x"ad",x"b7"),
   703 => (x"66",x"cc",x"87",x"ee"),
   704 => (x"f3",x"8e",x"ec",x"48"),
   705 => (x"5e",x"0e",x"87",x"d3"),
   706 => (x"0e",x"5d",x"5c",x"5b"),
   707 => (x"4b",x"71",x"86",x"f0"),
   708 => (x"4c",x"66",x"e0",x"c0"),
   709 => (x"9b",x"73",x"2c",x"c9"),
   710 => (x"87",x"e1",x"c3",x"02"),
   711 => (x"69",x"49",x"a3",x"c8"),
   712 => (x"87",x"d9",x"c3",x"02"),
   713 => (x"c0",x"49",x"a3",x"d0"),
   714 => (x"6b",x"79",x"66",x"e0"),
   715 => (x"c3",x"02",x"ac",x"7e"),
   716 => (x"c2",x"c3",x"87",x"cb"),
   717 => (x"ff",x"49",x"bf",x"ca"),
   718 => (x"74",x"4a",x"71",x"b9"),
   719 => (x"6e",x"48",x"71",x"9a"),
   720 => (x"58",x"a6",x"cc",x"98"),
   721 => (x"c4",x"4d",x"a3",x"c4"),
   722 => (x"78",x"6d",x"48",x"a6"),
   723 => (x"05",x"aa",x"66",x"c8"),
   724 => (x"7b",x"74",x"87",x"c5"),
   725 => (x"72",x"87",x"d1",x"c2"),
   726 => (x"fb",x"49",x"73",x"1e"),
   727 => (x"86",x"c4",x"87",x"e9"),
   728 => (x"c0",x"48",x"7e",x"70"),
   729 => (x"d0",x"04",x"a8",x"b7"),
   730 => (x"4a",x"a3",x"d4",x"87"),
   731 => (x"91",x"c8",x"49",x"6e"),
   732 => (x"21",x"49",x"a1",x"72"),
   733 => (x"c7",x"7d",x"69",x"7b"),
   734 => (x"cc",x"7b",x"c0",x"87"),
   735 => (x"7d",x"69",x"49",x"a3"),
   736 => (x"73",x"1e",x"66",x"c8"),
   737 => (x"87",x"ff",x"fa",x"49"),
   738 => (x"7e",x"70",x"86",x"c4"),
   739 => (x"49",x"a3",x"d4",x"c2"),
   740 => (x"69",x"48",x"a6",x"cc"),
   741 => (x"48",x"66",x"c8",x"78"),
   742 => (x"06",x"a8",x"66",x"cc"),
   743 => (x"48",x"6e",x"87",x"c9"),
   744 => (x"04",x"a8",x"b7",x"c0"),
   745 => (x"6e",x"87",x"e0",x"c0"),
   746 => (x"a8",x"b7",x"c0",x"48"),
   747 => (x"87",x"ec",x"c0",x"04"),
   748 => (x"6e",x"4a",x"a3",x"d4"),
   749 => (x"72",x"91",x"c8",x"49"),
   750 => (x"66",x"c8",x"49",x"a1"),
   751 => (x"70",x"88",x"69",x"48"),
   752 => (x"a9",x"66",x"cc",x"49"),
   753 => (x"73",x"87",x"d5",x"06"),
   754 => (x"87",x"c5",x"fb",x"49"),
   755 => (x"a3",x"d4",x"49",x"70"),
   756 => (x"72",x"91",x"c8",x"4a"),
   757 => (x"66",x"c8",x"49",x"a1"),
   758 => (x"79",x"66",x"c4",x"41"),
   759 => (x"49",x"74",x"8c",x"6b"),
   760 => (x"f5",x"49",x"73",x"1e"),
   761 => (x"86",x"c4",x"87",x"fa"),
   762 => (x"49",x"66",x"e0",x"c0"),
   763 => (x"02",x"99",x"ff",x"c7"),
   764 => (x"fa",x"c2",x"87",x"cb"),
   765 => (x"49",x"73",x"1e",x"c6"),
   766 => (x"c4",x"87",x"c6",x"f7"),
   767 => (x"ef",x"8e",x"f0",x"86"),
   768 => (x"73",x"1e",x"87",x"d7"),
   769 => (x"9b",x"4b",x"71",x"1e"),
   770 => (x"87",x"e4",x"c0",x"02"),
   771 => (x"5b",x"f3",x"c6",x"c3"),
   772 => (x"8a",x"c2",x"4a",x"73"),
   773 => (x"bf",x"c6",x"c2",x"c3"),
   774 => (x"c6",x"c3",x"92",x"49"),
   775 => (x"72",x"48",x"bf",x"df"),
   776 => (x"f7",x"c6",x"c3",x"80"),
   777 => (x"c4",x"48",x"71",x"58"),
   778 => (x"d6",x"c2",x"c3",x"30"),
   779 => (x"87",x"ed",x"c0",x"58"),
   780 => (x"48",x"ef",x"c6",x"c3"),
   781 => (x"bf",x"e3",x"c6",x"c3"),
   782 => (x"f3",x"c6",x"c3",x"78"),
   783 => (x"e7",x"c6",x"c3",x"48"),
   784 => (x"c2",x"c3",x"78",x"bf"),
   785 => (x"c9",x"02",x"bf",x"ce"),
   786 => (x"c6",x"c2",x"c3",x"87"),
   787 => (x"31",x"c4",x"49",x"bf"),
   788 => (x"c6",x"c3",x"87",x"c7"),
   789 => (x"c4",x"49",x"bf",x"eb"),
   790 => (x"d6",x"c2",x"c3",x"31"),
   791 => (x"87",x"fd",x"ed",x"59"),
   792 => (x"5c",x"5b",x"5e",x"0e"),
   793 => (x"c0",x"4a",x"71",x"0e"),
   794 => (x"02",x"9a",x"72",x"4b"),
   795 => (x"da",x"87",x"e1",x"c0"),
   796 => (x"69",x"9f",x"49",x"a2"),
   797 => (x"ce",x"c2",x"c3",x"4b"),
   798 => (x"87",x"cf",x"02",x"bf"),
   799 => (x"9f",x"49",x"a2",x"d4"),
   800 => (x"c0",x"4c",x"49",x"69"),
   801 => (x"d0",x"9c",x"ff",x"ff"),
   802 => (x"c0",x"87",x"c2",x"34"),
   803 => (x"b3",x"49",x"74",x"4c"),
   804 => (x"ed",x"fd",x"49",x"73"),
   805 => (x"87",x"c3",x"ed",x"87"),
   806 => (x"5c",x"5b",x"5e",x"0e"),
   807 => (x"86",x"f4",x"0e",x"5d"),
   808 => (x"7e",x"c0",x"4a",x"71"),
   809 => (x"d8",x"02",x"9a",x"72"),
   810 => (x"c2",x"fa",x"c2",x"87"),
   811 => (x"c2",x"78",x"c0",x"48"),
   812 => (x"c3",x"48",x"fa",x"f9"),
   813 => (x"78",x"bf",x"f3",x"c6"),
   814 => (x"48",x"fe",x"f9",x"c2"),
   815 => (x"bf",x"ef",x"c6",x"c3"),
   816 => (x"e3",x"c2",x"c3",x"78"),
   817 => (x"c3",x"50",x"c0",x"48"),
   818 => (x"49",x"bf",x"d2",x"c2"),
   819 => (x"bf",x"c2",x"fa",x"c2"),
   820 => (x"03",x"aa",x"71",x"4a"),
   821 => (x"72",x"87",x"c0",x"c4"),
   822 => (x"05",x"99",x"cf",x"49"),
   823 => (x"c2",x"87",x"e1",x"c0"),
   824 => (x"c2",x"1e",x"c6",x"fa"),
   825 => (x"49",x"bf",x"fa",x"f9"),
   826 => (x"48",x"fa",x"f9",x"c2"),
   827 => (x"71",x"78",x"a1",x"c1"),
   828 => (x"87",x"e7",x"dd",x"ff"),
   829 => (x"f9",x"c0",x"86",x"c4"),
   830 => (x"fa",x"c2",x"48",x"ec"),
   831 => (x"87",x"cc",x"78",x"c6"),
   832 => (x"bf",x"ec",x"f9",x"c0"),
   833 => (x"80",x"e0",x"c0",x"48"),
   834 => (x"58",x"f0",x"f9",x"c0"),
   835 => (x"bf",x"c2",x"fa",x"c2"),
   836 => (x"c2",x"80",x"c1",x"48"),
   837 => (x"27",x"58",x"c6",x"fa"),
   838 => (x"00",x"00",x"0e",x"6c"),
   839 => (x"4d",x"bf",x"97",x"bf"),
   840 => (x"e2",x"c2",x"02",x"9d"),
   841 => (x"ad",x"e5",x"c3",x"87"),
   842 => (x"87",x"db",x"c2",x"02"),
   843 => (x"bf",x"ec",x"f9",x"c0"),
   844 => (x"49",x"a3",x"cb",x"4b"),
   845 => (x"ac",x"cf",x"4c",x"11"),
   846 => (x"87",x"d2",x"c1",x"05"),
   847 => (x"99",x"df",x"49",x"75"),
   848 => (x"91",x"cd",x"89",x"c1"),
   849 => (x"81",x"d6",x"c2",x"c3"),
   850 => (x"12",x"4a",x"a3",x"c1"),
   851 => (x"4a",x"a3",x"c3",x"51"),
   852 => (x"a3",x"c5",x"51",x"12"),
   853 => (x"c7",x"51",x"12",x"4a"),
   854 => (x"51",x"12",x"4a",x"a3"),
   855 => (x"12",x"4a",x"a3",x"c9"),
   856 => (x"4a",x"a3",x"ce",x"51"),
   857 => (x"a3",x"d0",x"51",x"12"),
   858 => (x"d2",x"51",x"12",x"4a"),
   859 => (x"51",x"12",x"4a",x"a3"),
   860 => (x"12",x"4a",x"a3",x"d4"),
   861 => (x"4a",x"a3",x"d6",x"51"),
   862 => (x"a3",x"d8",x"51",x"12"),
   863 => (x"dc",x"51",x"12",x"4a"),
   864 => (x"51",x"12",x"4a",x"a3"),
   865 => (x"12",x"4a",x"a3",x"de"),
   866 => (x"c0",x"7e",x"c1",x"51"),
   867 => (x"49",x"74",x"87",x"f9"),
   868 => (x"c0",x"05",x"99",x"c8"),
   869 => (x"49",x"74",x"87",x"ea"),
   870 => (x"d0",x"05",x"99",x"d0"),
   871 => (x"02",x"66",x"dc",x"87"),
   872 => (x"73",x"87",x"ca",x"c0"),
   873 => (x"0f",x"66",x"dc",x"49"),
   874 => (x"d3",x"02",x"98",x"70"),
   875 => (x"c0",x"05",x"6e",x"87"),
   876 => (x"c2",x"c3",x"87",x"c6"),
   877 => (x"50",x"c0",x"48",x"d6"),
   878 => (x"bf",x"ec",x"f9",x"c0"),
   879 => (x"87",x"e7",x"c2",x"48"),
   880 => (x"48",x"e3",x"c2",x"c3"),
   881 => (x"c3",x"7e",x"50",x"c0"),
   882 => (x"49",x"bf",x"d2",x"c2"),
   883 => (x"bf",x"c2",x"fa",x"c2"),
   884 => (x"04",x"aa",x"71",x"4a"),
   885 => (x"c3",x"87",x"c0",x"fc"),
   886 => (x"05",x"bf",x"f3",x"c6"),
   887 => (x"c3",x"87",x"c8",x"c0"),
   888 => (x"02",x"bf",x"ce",x"c2"),
   889 => (x"c0",x"87",x"fe",x"c1"),
   890 => (x"ff",x"48",x"f0",x"f9"),
   891 => (x"fe",x"f9",x"c2",x"78"),
   892 => (x"ec",x"e7",x"49",x"bf"),
   893 => (x"c2",x"49",x"70",x"87"),
   894 => (x"c4",x"59",x"c2",x"fa"),
   895 => (x"f9",x"c2",x"48",x"a6"),
   896 => (x"c3",x"78",x"bf",x"fe"),
   897 => (x"02",x"bf",x"ce",x"c2"),
   898 => (x"c4",x"87",x"d8",x"c0"),
   899 => (x"ff",x"cf",x"49",x"66"),
   900 => (x"99",x"f8",x"ff",x"ff"),
   901 => (x"c5",x"c0",x"02",x"a9"),
   902 => (x"c0",x"4d",x"c0",x"87"),
   903 => (x"4d",x"c1",x"87",x"e1"),
   904 => (x"c4",x"87",x"dc",x"c0"),
   905 => (x"ff",x"cf",x"49",x"66"),
   906 => (x"02",x"a9",x"99",x"f8"),
   907 => (x"c8",x"87",x"c8",x"c0"),
   908 => (x"78",x"c0",x"48",x"a6"),
   909 => (x"c8",x"87",x"c5",x"c0"),
   910 => (x"78",x"c1",x"48",x"a6"),
   911 => (x"75",x"4d",x"66",x"c8"),
   912 => (x"e0",x"c0",x"05",x"9d"),
   913 => (x"49",x"66",x"c4",x"87"),
   914 => (x"c2",x"c3",x"89",x"c2"),
   915 => (x"91",x"4a",x"bf",x"c6"),
   916 => (x"bf",x"df",x"c6",x"c3"),
   917 => (x"fa",x"f9",x"c2",x"4a"),
   918 => (x"78",x"a1",x"72",x"48"),
   919 => (x"48",x"c2",x"fa",x"c2"),
   920 => (x"e2",x"f9",x"78",x"c0"),
   921 => (x"f4",x"48",x"c0",x"87"),
   922 => (x"87",x"ed",x"e5",x"8e"),
   923 => (x"00",x"00",x"00",x"00"),
   924 => (x"ff",x"ff",x"ff",x"ff"),
   925 => (x"00",x"00",x"0e",x"7c"),
   926 => (x"00",x"00",x"0e",x"85"),
   927 => (x"33",x"54",x"41",x"46"),
   928 => (x"20",x"20",x"20",x"32"),
   929 => (x"54",x"41",x"46",x"00"),
   930 => (x"20",x"20",x"36",x"31"),
   931 => (x"ff",x"1e",x"00",x"20"),
   932 => (x"ff",x"c3",x"48",x"d4"),
   933 => (x"26",x"48",x"68",x"78"),
   934 => (x"d4",x"ff",x"1e",x"4f"),
   935 => (x"78",x"ff",x"c3",x"48"),
   936 => (x"c8",x"48",x"d0",x"ff"),
   937 => (x"d4",x"ff",x"78",x"e1"),
   938 => (x"c3",x"78",x"d4",x"48"),
   939 => (x"ff",x"48",x"f7",x"c6"),
   940 => (x"26",x"50",x"bf",x"d4"),
   941 => (x"d0",x"ff",x"1e",x"4f"),
   942 => (x"78",x"e0",x"c0",x"48"),
   943 => (x"ff",x"1e",x"4f",x"26"),
   944 => (x"49",x"70",x"87",x"cc"),
   945 => (x"87",x"c6",x"02",x"99"),
   946 => (x"05",x"a9",x"fb",x"c0"),
   947 => (x"48",x"71",x"87",x"f1"),
   948 => (x"5e",x"0e",x"4f",x"26"),
   949 => (x"71",x"0e",x"5c",x"5b"),
   950 => (x"fe",x"4c",x"c0",x"4b"),
   951 => (x"49",x"70",x"87",x"f0"),
   952 => (x"f9",x"c0",x"02",x"99"),
   953 => (x"a9",x"ec",x"c0",x"87"),
   954 => (x"87",x"f2",x"c0",x"02"),
   955 => (x"02",x"a9",x"fb",x"c0"),
   956 => (x"cc",x"87",x"eb",x"c0"),
   957 => (x"03",x"ac",x"b7",x"66"),
   958 => (x"66",x"d0",x"87",x"c7"),
   959 => (x"71",x"87",x"c2",x"02"),
   960 => (x"02",x"99",x"71",x"53"),
   961 => (x"84",x"c1",x"87",x"c2"),
   962 => (x"70",x"87",x"c3",x"fe"),
   963 => (x"cd",x"02",x"99",x"49"),
   964 => (x"a9",x"ec",x"c0",x"87"),
   965 => (x"c0",x"87",x"c7",x"02"),
   966 => (x"ff",x"05",x"a9",x"fb"),
   967 => (x"66",x"d0",x"87",x"d5"),
   968 => (x"c0",x"87",x"c3",x"02"),
   969 => (x"ec",x"c0",x"7b",x"97"),
   970 => (x"87",x"c4",x"05",x"a9"),
   971 => (x"87",x"c5",x"4a",x"74"),
   972 => (x"0a",x"c0",x"4a",x"74"),
   973 => (x"c2",x"48",x"72",x"8a"),
   974 => (x"26",x"4d",x"26",x"87"),
   975 => (x"26",x"4b",x"26",x"4c"),
   976 => (x"c9",x"fd",x"1e",x"4f"),
   977 => (x"c0",x"49",x"70",x"87"),
   978 => (x"04",x"a9",x"b7",x"f0"),
   979 => (x"f9",x"c0",x"87",x"ca"),
   980 => (x"c3",x"01",x"a9",x"b7"),
   981 => (x"89",x"f0",x"c0",x"87"),
   982 => (x"a9",x"b7",x"c1",x"c1"),
   983 => (x"c1",x"87",x"ca",x"04"),
   984 => (x"01",x"a9",x"b7",x"da"),
   985 => (x"f7",x"c0",x"87",x"c3"),
   986 => (x"26",x"48",x"71",x"89"),
   987 => (x"5b",x"5e",x"0e",x"4f"),
   988 => (x"4a",x"71",x"0e",x"5c"),
   989 => (x"72",x"4c",x"d4",x"ff"),
   990 => (x"87",x"ea",x"c0",x"49"),
   991 => (x"02",x"9b",x"4b",x"70"),
   992 => (x"8b",x"c1",x"87",x"c2"),
   993 => (x"c8",x"48",x"d0",x"ff"),
   994 => (x"d5",x"c1",x"78",x"c5"),
   995 => (x"c6",x"49",x"73",x"7c"),
   996 => (x"c5",x"e2",x"c2",x"31"),
   997 => (x"48",x"4a",x"bf",x"97"),
   998 => (x"7c",x"70",x"b0",x"71"),
   999 => (x"c4",x"48",x"d0",x"ff"),
  1000 => (x"fe",x"48",x"73",x"78"),
  1001 => (x"5e",x"0e",x"87",x"d5"),
  1002 => (x"0e",x"5d",x"5c",x"5b"),
  1003 => (x"4c",x"71",x"86",x"f8"),
  1004 => (x"e4",x"fb",x"7e",x"c0"),
  1005 => (x"c1",x"4b",x"c0",x"87"),
  1006 => (x"bf",x"97",x"d3",x"c1"),
  1007 => (x"04",x"a9",x"c0",x"49"),
  1008 => (x"f9",x"fb",x"87",x"cf"),
  1009 => (x"c1",x"83",x"c1",x"87"),
  1010 => (x"bf",x"97",x"d3",x"c1"),
  1011 => (x"f1",x"06",x"ab",x"49"),
  1012 => (x"d3",x"c1",x"c1",x"87"),
  1013 => (x"cf",x"02",x"bf",x"97"),
  1014 => (x"87",x"f2",x"fa",x"87"),
  1015 => (x"02",x"99",x"49",x"70"),
  1016 => (x"ec",x"c0",x"87",x"c6"),
  1017 => (x"87",x"f1",x"05",x"a9"),
  1018 => (x"e1",x"fa",x"4b",x"c0"),
  1019 => (x"fa",x"4d",x"70",x"87"),
  1020 => (x"a6",x"c8",x"87",x"dc"),
  1021 => (x"87",x"d6",x"fa",x"58"),
  1022 => (x"83",x"c1",x"4a",x"70"),
  1023 => (x"97",x"49",x"a4",x"c8"),
  1024 => (x"02",x"ad",x"49",x"69"),
  1025 => (x"ff",x"c0",x"87",x"c7"),
  1026 => (x"e7",x"c0",x"05",x"ad"),
  1027 => (x"49",x"a4",x"c9",x"87"),
  1028 => (x"c4",x"49",x"69",x"97"),
  1029 => (x"c7",x"02",x"a9",x"66"),
  1030 => (x"ff",x"c0",x"48",x"87"),
  1031 => (x"87",x"d4",x"05",x"a8"),
  1032 => (x"97",x"49",x"a4",x"ca"),
  1033 => (x"02",x"aa",x"49",x"69"),
  1034 => (x"ff",x"c0",x"87",x"c6"),
  1035 => (x"87",x"c4",x"05",x"aa"),
  1036 => (x"87",x"d0",x"7e",x"c1"),
  1037 => (x"02",x"ad",x"ec",x"c0"),
  1038 => (x"fb",x"c0",x"87",x"c6"),
  1039 => (x"87",x"c4",x"05",x"ad"),
  1040 => (x"7e",x"c1",x"4b",x"c0"),
  1041 => (x"e1",x"fe",x"02",x"6e"),
  1042 => (x"87",x"e9",x"f9",x"87"),
  1043 => (x"8e",x"f8",x"48",x"73"),
  1044 => (x"00",x"87",x"e6",x"fb"),
  1045 => (x"5c",x"5b",x"5e",x"0e"),
  1046 => (x"71",x"1e",x"0e",x"5d"),
  1047 => (x"4d",x"4c",x"c0",x"4b"),
  1048 => (x"e8",x"c0",x"04",x"ab"),
  1049 => (x"e6",x"fe",x"c0",x"87"),
  1050 => (x"02",x"9d",x"75",x"1e"),
  1051 => (x"4a",x"c0",x"87",x"c4"),
  1052 => (x"4a",x"c1",x"87",x"c2"),
  1053 => (x"df",x"f0",x"49",x"72"),
  1054 => (x"70",x"86",x"c4",x"87"),
  1055 => (x"6e",x"84",x"c1",x"7e"),
  1056 => (x"73",x"87",x"c2",x"05"),
  1057 => (x"73",x"85",x"c1",x"4c"),
  1058 => (x"d8",x"ff",x"06",x"ac"),
  1059 => (x"26",x"48",x"6e",x"87"),
  1060 => (x"4c",x"26",x"4d",x"26"),
  1061 => (x"4f",x"26",x"4b",x"26"),
  1062 => (x"5c",x"5b",x"5e",x"0e"),
  1063 => (x"71",x"1e",x"0e",x"5d"),
  1064 => (x"91",x"de",x"49",x"4c"),
  1065 => (x"4d",x"d1",x"c7",x"c3"),
  1066 => (x"6d",x"97",x"85",x"71"),
  1067 => (x"87",x"dd",x"c1",x"02"),
  1068 => (x"bf",x"fc",x"c6",x"c3"),
  1069 => (x"72",x"82",x"74",x"4a"),
  1070 => (x"87",x"d8",x"fe",x"49"),
  1071 => (x"02",x"6e",x"7e",x"70"),
  1072 => (x"c3",x"87",x"f3",x"c0"),
  1073 => (x"6e",x"4b",x"c4",x"c7"),
  1074 => (x"fe",x"49",x"cb",x"4a"),
  1075 => (x"74",x"87",x"d9",x"ff"),
  1076 => (x"c1",x"93",x"cb",x"4b"),
  1077 => (x"c4",x"83",x"dc",x"e4"),
  1078 => (x"d1",x"c4",x"c1",x"83"),
  1079 => (x"c1",x"49",x"74",x"7b"),
  1080 => (x"75",x"87",x"fe",x"c2"),
  1081 => (x"d0",x"c7",x"c3",x"7b"),
  1082 => (x"1e",x"49",x"bf",x"97"),
  1083 => (x"49",x"c4",x"c7",x"c3"),
  1084 => (x"87",x"d3",x"dd",x"c1"),
  1085 => (x"49",x"74",x"86",x"c4"),
  1086 => (x"87",x"e5",x"c2",x"c1"),
  1087 => (x"c4",x"c1",x"49",x"c0"),
  1088 => (x"c6",x"c3",x"87",x"c4"),
  1089 => (x"78",x"c0",x"48",x"f8"),
  1090 => (x"fa",x"dc",x"49",x"c1"),
  1091 => (x"ff",x"fd",x"26",x"87"),
  1092 => (x"61",x"6f",x"4c",x"87"),
  1093 => (x"67",x"6e",x"69",x"64"),
  1094 => (x"00",x"2e",x"2e",x"2e"),
  1095 => (x"5c",x"5b",x"5e",x"0e"),
  1096 => (x"4a",x"4b",x"71",x"0e"),
  1097 => (x"bf",x"fc",x"c6",x"c3"),
  1098 => (x"fc",x"49",x"72",x"82"),
  1099 => (x"4c",x"70",x"87",x"e6"),
  1100 => (x"87",x"c4",x"02",x"9c"),
  1101 => (x"87",x"e8",x"ec",x"49"),
  1102 => (x"48",x"fc",x"c6",x"c3"),
  1103 => (x"49",x"c1",x"78",x"c0"),
  1104 => (x"fd",x"87",x"c4",x"dc"),
  1105 => (x"5e",x"0e",x"87",x"cc"),
  1106 => (x"0e",x"5d",x"5c",x"5b"),
  1107 => (x"fa",x"c2",x"86",x"f4"),
  1108 => (x"4c",x"c0",x"4d",x"c6"),
  1109 => (x"c0",x"48",x"a6",x"c4"),
  1110 => (x"fc",x"c6",x"c3",x"78"),
  1111 => (x"a9",x"c0",x"49",x"bf"),
  1112 => (x"87",x"c1",x"c1",x"06"),
  1113 => (x"48",x"c6",x"fa",x"c2"),
  1114 => (x"f8",x"c0",x"02",x"98"),
  1115 => (x"e6",x"fe",x"c0",x"87"),
  1116 => (x"02",x"66",x"c8",x"1e"),
  1117 => (x"a6",x"c4",x"87",x"c7"),
  1118 => (x"c5",x"78",x"c0",x"48"),
  1119 => (x"48",x"a6",x"c4",x"87"),
  1120 => (x"66",x"c4",x"78",x"c1"),
  1121 => (x"87",x"d0",x"ec",x"49"),
  1122 => (x"4d",x"70",x"86",x"c4"),
  1123 => (x"66",x"c4",x"84",x"c1"),
  1124 => (x"c8",x"80",x"c1",x"48"),
  1125 => (x"c6",x"c3",x"58",x"a6"),
  1126 => (x"ac",x"49",x"bf",x"fc"),
  1127 => (x"75",x"87",x"c6",x"03"),
  1128 => (x"c8",x"ff",x"05",x"9d"),
  1129 => (x"75",x"4c",x"c0",x"87"),
  1130 => (x"e0",x"c3",x"02",x"9d"),
  1131 => (x"e6",x"fe",x"c0",x"87"),
  1132 => (x"02",x"66",x"c8",x"1e"),
  1133 => (x"a6",x"cc",x"87",x"c7"),
  1134 => (x"c5",x"78",x"c0",x"48"),
  1135 => (x"48",x"a6",x"cc",x"87"),
  1136 => (x"66",x"cc",x"78",x"c1"),
  1137 => (x"87",x"d0",x"eb",x"49"),
  1138 => (x"7e",x"70",x"86",x"c4"),
  1139 => (x"e9",x"c2",x"02",x"6e"),
  1140 => (x"cb",x"49",x"6e",x"87"),
  1141 => (x"49",x"69",x"97",x"81"),
  1142 => (x"c1",x"02",x"99",x"d0"),
  1143 => (x"c4",x"c1",x"87",x"d6"),
  1144 => (x"49",x"74",x"4a",x"dc"),
  1145 => (x"e4",x"c1",x"91",x"cb"),
  1146 => (x"79",x"72",x"81",x"dc"),
  1147 => (x"ff",x"c3",x"81",x"c8"),
  1148 => (x"de",x"49",x"74",x"51"),
  1149 => (x"d1",x"c7",x"c3",x"91"),
  1150 => (x"c2",x"85",x"71",x"4d"),
  1151 => (x"c1",x"7d",x"97",x"c1"),
  1152 => (x"e0",x"c0",x"49",x"a5"),
  1153 => (x"d6",x"c2",x"c3",x"51"),
  1154 => (x"d2",x"02",x"bf",x"97"),
  1155 => (x"c2",x"84",x"c1",x"87"),
  1156 => (x"c2",x"c3",x"4b",x"a5"),
  1157 => (x"49",x"db",x"4a",x"d6"),
  1158 => (x"87",x"cc",x"fa",x"fe"),
  1159 => (x"cd",x"87",x"db",x"c1"),
  1160 => (x"51",x"c0",x"49",x"a5"),
  1161 => (x"a5",x"c2",x"84",x"c1"),
  1162 => (x"cb",x"4a",x"6e",x"4b"),
  1163 => (x"f7",x"f9",x"fe",x"49"),
  1164 => (x"87",x"c6",x"c1",x"87"),
  1165 => (x"4a",x"d8",x"c2",x"c1"),
  1166 => (x"91",x"cb",x"49",x"74"),
  1167 => (x"81",x"dc",x"e4",x"c1"),
  1168 => (x"c2",x"c3",x"79",x"72"),
  1169 => (x"02",x"bf",x"97",x"d6"),
  1170 => (x"49",x"74",x"87",x"d8"),
  1171 => (x"84",x"c1",x"91",x"de"),
  1172 => (x"4b",x"d1",x"c7",x"c3"),
  1173 => (x"c2",x"c3",x"83",x"71"),
  1174 => (x"49",x"dd",x"4a",x"d6"),
  1175 => (x"87",x"c8",x"f9",x"fe"),
  1176 => (x"4b",x"74",x"87",x"d8"),
  1177 => (x"c7",x"c3",x"93",x"de"),
  1178 => (x"a3",x"cb",x"83",x"d1"),
  1179 => (x"c1",x"51",x"c0",x"49"),
  1180 => (x"4a",x"6e",x"73",x"84"),
  1181 => (x"f8",x"fe",x"49",x"cb"),
  1182 => (x"66",x"c4",x"87",x"ee"),
  1183 => (x"c8",x"80",x"c1",x"48"),
  1184 => (x"ac",x"c7",x"58",x"a6"),
  1185 => (x"87",x"c5",x"c0",x"03"),
  1186 => (x"e0",x"fc",x"05",x"6e"),
  1187 => (x"f4",x"48",x"74",x"87"),
  1188 => (x"87",x"fc",x"f7",x"8e"),
  1189 => (x"71",x"1e",x"73",x"1e"),
  1190 => (x"91",x"cb",x"49",x"4b"),
  1191 => (x"81",x"dc",x"e4",x"c1"),
  1192 => (x"c2",x"4a",x"a1",x"c8"),
  1193 => (x"12",x"48",x"c5",x"e2"),
  1194 => (x"4a",x"a1",x"c9",x"50"),
  1195 => (x"48",x"d3",x"c1",x"c1"),
  1196 => (x"81",x"ca",x"50",x"12"),
  1197 => (x"48",x"d0",x"c7",x"c3"),
  1198 => (x"c7",x"c3",x"50",x"11"),
  1199 => (x"49",x"bf",x"97",x"d0"),
  1200 => (x"c1",x"49",x"c0",x"1e"),
  1201 => (x"c3",x"87",x"c0",x"d6"),
  1202 => (x"de",x"48",x"f8",x"c6"),
  1203 => (x"d5",x"49",x"c1",x"78"),
  1204 => (x"f6",x"26",x"87",x"f5"),
  1205 => (x"71",x"1e",x"87",x"fe"),
  1206 => (x"91",x"cb",x"49",x"4a"),
  1207 => (x"81",x"dc",x"e4",x"c1"),
  1208 => (x"48",x"11",x"81",x"c8"),
  1209 => (x"58",x"fc",x"c6",x"c3"),
  1210 => (x"48",x"fc",x"c6",x"c3"),
  1211 => (x"49",x"c1",x"78",x"c0"),
  1212 => (x"26",x"87",x"d4",x"d5"),
  1213 => (x"49",x"c0",x"1e",x"4f"),
  1214 => (x"87",x"ca",x"fc",x"c0"),
  1215 => (x"71",x"1e",x"4f",x"26"),
  1216 => (x"87",x"d2",x"02",x"99"),
  1217 => (x"48",x"f1",x"e5",x"c1"),
  1218 => (x"80",x"f7",x"50",x"c0"),
  1219 => (x"40",x"d6",x"cb",x"c1"),
  1220 => (x"78",x"d5",x"e4",x"c1"),
  1221 => (x"e5",x"c1",x"87",x"ce"),
  1222 => (x"e4",x"c1",x"48",x"ed"),
  1223 => (x"80",x"fc",x"78",x"ce"),
  1224 => (x"78",x"f5",x"cb",x"c1"),
  1225 => (x"5e",x"0e",x"4f",x"26"),
  1226 => (x"71",x"0e",x"5c",x"5b"),
  1227 => (x"92",x"cb",x"4a",x"4c"),
  1228 => (x"82",x"dc",x"e4",x"c1"),
  1229 => (x"c9",x"49",x"a2",x"c8"),
  1230 => (x"6b",x"97",x"4b",x"a2"),
  1231 => (x"69",x"97",x"1e",x"4b"),
  1232 => (x"82",x"ca",x"1e",x"49"),
  1233 => (x"e7",x"c0",x"49",x"12"),
  1234 => (x"49",x"c0",x"87",x"c5"),
  1235 => (x"74",x"87",x"f8",x"d3"),
  1236 => (x"cc",x"f9",x"c0",x"49"),
  1237 => (x"f4",x"8e",x"f8",x"87"),
  1238 => (x"73",x"1e",x"87",x"f8"),
  1239 => (x"c6",x"4b",x"71",x"1e"),
  1240 => (x"db",x"02",x"4a",x"a3"),
  1241 => (x"02",x"8a",x"c1",x"87"),
  1242 => (x"02",x"8a",x"87",x"d6"),
  1243 => (x"8a",x"87",x"da",x"c1"),
  1244 => (x"87",x"fc",x"c0",x"02"),
  1245 => (x"e1",x"c0",x"02",x"8a"),
  1246 => (x"cb",x"02",x"8a",x"87"),
  1247 => (x"87",x"db",x"c1",x"87"),
  1248 => (x"d1",x"fd",x"49",x"c7"),
  1249 => (x"87",x"de",x"c1",x"87"),
  1250 => (x"bf",x"fc",x"c6",x"c3"),
  1251 => (x"87",x"cb",x"c1",x"02"),
  1252 => (x"c3",x"88",x"c1",x"48"),
  1253 => (x"c1",x"58",x"c0",x"c7"),
  1254 => (x"c7",x"c3",x"87",x"c1"),
  1255 => (x"c0",x"02",x"bf",x"c0"),
  1256 => (x"c6",x"c3",x"87",x"f9"),
  1257 => (x"c1",x"48",x"bf",x"fc"),
  1258 => (x"c0",x"c7",x"c3",x"80"),
  1259 => (x"87",x"eb",x"c0",x"58"),
  1260 => (x"bf",x"fc",x"c6",x"c3"),
  1261 => (x"c3",x"89",x"c6",x"49"),
  1262 => (x"c0",x"59",x"c0",x"c7"),
  1263 => (x"da",x"03",x"a9",x"b7"),
  1264 => (x"fc",x"c6",x"c3",x"87"),
  1265 => (x"d2",x"78",x"c0",x"48"),
  1266 => (x"c0",x"c7",x"c3",x"87"),
  1267 => (x"87",x"cb",x"02",x"bf"),
  1268 => (x"bf",x"fc",x"c6",x"c3"),
  1269 => (x"c3",x"80",x"c6",x"48"),
  1270 => (x"c0",x"58",x"c0",x"c7"),
  1271 => (x"87",x"e7",x"d1",x"49"),
  1272 => (x"f6",x"c0",x"49",x"73"),
  1273 => (x"eb",x"f2",x"87",x"fb"),
  1274 => (x"5b",x"5e",x"0e",x"87"),
  1275 => (x"4c",x"71",x"0e",x"5c"),
  1276 => (x"74",x"1e",x"66",x"cc"),
  1277 => (x"c1",x"93",x"cb",x"4b"),
  1278 => (x"c4",x"83",x"dc",x"e4"),
  1279 => (x"49",x"6a",x"4a",x"a3"),
  1280 => (x"87",x"f4",x"f2",x"fe"),
  1281 => (x"7b",x"d4",x"ca",x"c1"),
  1282 => (x"d4",x"49",x"a3",x"c8"),
  1283 => (x"a3",x"c9",x"51",x"66"),
  1284 => (x"51",x"66",x"d8",x"49"),
  1285 => (x"dc",x"49",x"a3",x"ca"),
  1286 => (x"f1",x"26",x"51",x"66"),
  1287 => (x"5e",x"0e",x"87",x"f4"),
  1288 => (x"0e",x"5d",x"5c",x"5b"),
  1289 => (x"d8",x"86",x"d0",x"ff"),
  1290 => (x"a6",x"c4",x"59",x"a6"),
  1291 => (x"c4",x"78",x"c0",x"48"),
  1292 => (x"66",x"c4",x"c1",x"80"),
  1293 => (x"c1",x"80",x"c4",x"78"),
  1294 => (x"c1",x"80",x"c4",x"78"),
  1295 => (x"c0",x"c7",x"c3",x"78"),
  1296 => (x"c3",x"78",x"c1",x"48"),
  1297 => (x"48",x"bf",x"f8",x"c6"),
  1298 => (x"cb",x"05",x"a8",x"de"),
  1299 => (x"87",x"f6",x"f3",x"87"),
  1300 => (x"a6",x"c8",x"49",x"70"),
  1301 => (x"87",x"f8",x"ce",x"59"),
  1302 => (x"e9",x"87",x"fe",x"e8"),
  1303 => (x"ed",x"e8",x"87",x"e0"),
  1304 => (x"c0",x"4c",x"70",x"87"),
  1305 => (x"c1",x"02",x"ac",x"fb"),
  1306 => (x"66",x"d4",x"87",x"d0"),
  1307 => (x"87",x"c2",x"c1",x"05"),
  1308 => (x"c1",x"1e",x"1e",x"c0"),
  1309 => (x"ff",x"e5",x"c1",x"1e"),
  1310 => (x"fd",x"49",x"c0",x"1e"),
  1311 => (x"d0",x"c1",x"87",x"eb"),
  1312 => (x"82",x"c4",x"4a",x"66"),
  1313 => (x"81",x"c7",x"49",x"6a"),
  1314 => (x"1e",x"c1",x"51",x"74"),
  1315 => (x"49",x"6a",x"1e",x"d8"),
  1316 => (x"fd",x"e8",x"81",x"c8"),
  1317 => (x"c1",x"86",x"d8",x"87"),
  1318 => (x"c0",x"48",x"66",x"c4"),
  1319 => (x"87",x"c7",x"01",x"a8"),
  1320 => (x"c1",x"48",x"a6",x"c4"),
  1321 => (x"c1",x"87",x"ce",x"78"),
  1322 => (x"c1",x"48",x"66",x"c4"),
  1323 => (x"58",x"a6",x"cc",x"88"),
  1324 => (x"c9",x"e8",x"87",x"c3"),
  1325 => (x"48",x"a6",x"cc",x"87"),
  1326 => (x"9c",x"74",x"78",x"c2"),
  1327 => (x"87",x"cc",x"cd",x"02"),
  1328 => (x"c1",x"48",x"66",x"c4"),
  1329 => (x"03",x"a8",x"66",x"c8"),
  1330 => (x"d8",x"87",x"c1",x"cd"),
  1331 => (x"78",x"c0",x"48",x"a6"),
  1332 => (x"70",x"87",x"fb",x"e6"),
  1333 => (x"ac",x"d0",x"c1",x"4c"),
  1334 => (x"87",x"d6",x"c2",x"05"),
  1335 => (x"e9",x"7e",x"66",x"d8"),
  1336 => (x"49",x"70",x"87",x"df"),
  1337 => (x"e6",x"59",x"a6",x"dc"),
  1338 => (x"4c",x"70",x"87",x"e4"),
  1339 => (x"05",x"ac",x"ec",x"c0"),
  1340 => (x"c4",x"87",x"ea",x"c1"),
  1341 => (x"91",x"cb",x"49",x"66"),
  1342 => (x"81",x"66",x"c0",x"c1"),
  1343 => (x"6a",x"4a",x"a1",x"c4"),
  1344 => (x"4a",x"a1",x"c8",x"4d"),
  1345 => (x"c1",x"52",x"66",x"d8"),
  1346 => (x"e6",x"79",x"d6",x"cb"),
  1347 => (x"4c",x"70",x"87",x"c0"),
  1348 => (x"87",x"d8",x"02",x"9c"),
  1349 => (x"02",x"ac",x"fb",x"c0"),
  1350 => (x"55",x"74",x"87",x"d2"),
  1351 => (x"70",x"87",x"ef",x"e5"),
  1352 => (x"c7",x"02",x"9c",x"4c"),
  1353 => (x"ac",x"fb",x"c0",x"87"),
  1354 => (x"87",x"ee",x"ff",x"05"),
  1355 => (x"c2",x"55",x"e0",x"c0"),
  1356 => (x"97",x"c0",x"55",x"c1"),
  1357 => (x"49",x"66",x"d4",x"7d"),
  1358 => (x"db",x"05",x"a9",x"6e"),
  1359 => (x"48",x"66",x"c4",x"87"),
  1360 => (x"04",x"a8",x"66",x"c8"),
  1361 => (x"66",x"c4",x"87",x"ca"),
  1362 => (x"c8",x"80",x"c1",x"48"),
  1363 => (x"87",x"c8",x"58",x"a6"),
  1364 => (x"c1",x"48",x"66",x"c8"),
  1365 => (x"58",x"a6",x"cc",x"88"),
  1366 => (x"70",x"87",x"f3",x"e4"),
  1367 => (x"ac",x"d0",x"c1",x"4c"),
  1368 => (x"d0",x"87",x"c8",x"05"),
  1369 => (x"80",x"c1",x"48",x"66"),
  1370 => (x"c1",x"58",x"a6",x"d4"),
  1371 => (x"fd",x"02",x"ac",x"d0"),
  1372 => (x"a6",x"dc",x"87",x"ea"),
  1373 => (x"78",x"66",x"d4",x"48"),
  1374 => (x"dc",x"48",x"66",x"d8"),
  1375 => (x"c9",x"05",x"a8",x"66"),
  1376 => (x"e0",x"c0",x"87",x"dc"),
  1377 => (x"f0",x"c0",x"48",x"a6"),
  1378 => (x"cc",x"80",x"c4",x"78"),
  1379 => (x"80",x"c4",x"78",x"66"),
  1380 => (x"74",x"7e",x"78",x"c0"),
  1381 => (x"88",x"fb",x"c0",x"48"),
  1382 => (x"58",x"a6",x"f0",x"c0"),
  1383 => (x"c8",x"02",x"98",x"70"),
  1384 => (x"cb",x"48",x"87",x"d7"),
  1385 => (x"a6",x"f0",x"c0",x"88"),
  1386 => (x"02",x"98",x"70",x"58"),
  1387 => (x"48",x"87",x"e9",x"c0"),
  1388 => (x"f0",x"c0",x"88",x"c9"),
  1389 => (x"98",x"70",x"58",x"a6"),
  1390 => (x"87",x"e1",x"c3",x"02"),
  1391 => (x"c0",x"88",x"c4",x"48"),
  1392 => (x"70",x"58",x"a6",x"f0"),
  1393 => (x"87",x"de",x"02",x"98"),
  1394 => (x"c0",x"88",x"c1",x"48"),
  1395 => (x"70",x"58",x"a6",x"f0"),
  1396 => (x"c8",x"c3",x"02",x"98"),
  1397 => (x"87",x"db",x"c7",x"87"),
  1398 => (x"48",x"a6",x"e0",x"c0"),
  1399 => (x"66",x"cc",x"78",x"c0"),
  1400 => (x"d0",x"80",x"c1",x"48"),
  1401 => (x"e5",x"e2",x"58",x"a6"),
  1402 => (x"c0",x"4c",x"70",x"87"),
  1403 => (x"d5",x"02",x"ac",x"ec"),
  1404 => (x"66",x"e0",x"c0",x"87"),
  1405 => (x"c0",x"87",x"c6",x"02"),
  1406 => (x"c9",x"5c",x"a6",x"e4"),
  1407 => (x"c0",x"48",x"74",x"87"),
  1408 => (x"e8",x"c0",x"88",x"f0"),
  1409 => (x"ec",x"c0",x"58",x"a6"),
  1410 => (x"87",x"cc",x"02",x"ac"),
  1411 => (x"70",x"87",x"ff",x"e1"),
  1412 => (x"ac",x"ec",x"c0",x"4c"),
  1413 => (x"87",x"f4",x"ff",x"05"),
  1414 => (x"1e",x"66",x"e0",x"c0"),
  1415 => (x"1e",x"49",x"66",x"d4"),
  1416 => (x"1e",x"66",x"ec",x"c0"),
  1417 => (x"1e",x"ff",x"e5",x"c1"),
  1418 => (x"f6",x"49",x"66",x"d4"),
  1419 => (x"1e",x"c0",x"87",x"fb"),
  1420 => (x"66",x"dc",x"1e",x"ca"),
  1421 => (x"c1",x"91",x"cb",x"49"),
  1422 => (x"d8",x"81",x"66",x"d8"),
  1423 => (x"a1",x"c4",x"48",x"a6"),
  1424 => (x"bf",x"66",x"d8",x"78"),
  1425 => (x"87",x"ca",x"e2",x"49"),
  1426 => (x"b7",x"c0",x"86",x"d8"),
  1427 => (x"c7",x"c1",x"06",x"a8"),
  1428 => (x"de",x"1e",x"c1",x"87"),
  1429 => (x"bf",x"66",x"c8",x"1e"),
  1430 => (x"87",x"f6",x"e1",x"49"),
  1431 => (x"49",x"70",x"86",x"c8"),
  1432 => (x"88",x"08",x"c0",x"48"),
  1433 => (x"58",x"a6",x"e4",x"c0"),
  1434 => (x"06",x"a8",x"b7",x"c0"),
  1435 => (x"c0",x"87",x"e9",x"c0"),
  1436 => (x"dd",x"48",x"66",x"e0"),
  1437 => (x"df",x"03",x"a8",x"b7"),
  1438 => (x"49",x"bf",x"6e",x"87"),
  1439 => (x"81",x"66",x"e0",x"c0"),
  1440 => (x"66",x"51",x"e0",x"c0"),
  1441 => (x"6e",x"81",x"c1",x"49"),
  1442 => (x"c1",x"c2",x"81",x"bf"),
  1443 => (x"66",x"e0",x"c0",x"51"),
  1444 => (x"6e",x"81",x"c2",x"49"),
  1445 => (x"51",x"c0",x"81",x"bf"),
  1446 => (x"dc",x"c4",x"7e",x"c1"),
  1447 => (x"87",x"e1",x"e2",x"87"),
  1448 => (x"58",x"a6",x"e4",x"c0"),
  1449 => (x"c0",x"87",x"da",x"e2"),
  1450 => (x"c0",x"58",x"a6",x"e8"),
  1451 => (x"c0",x"05",x"a8",x"ec"),
  1452 => (x"e4",x"c0",x"87",x"cb"),
  1453 => (x"e0",x"c0",x"48",x"a6"),
  1454 => (x"c4",x"c0",x"78",x"66"),
  1455 => (x"cd",x"df",x"ff",x"87"),
  1456 => (x"49",x"66",x"c4",x"87"),
  1457 => (x"c0",x"c1",x"91",x"cb"),
  1458 => (x"80",x"71",x"48",x"66"),
  1459 => (x"4a",x"6e",x"7e",x"70"),
  1460 => (x"49",x"6e",x"82",x"c8"),
  1461 => (x"e0",x"c0",x"81",x"ca"),
  1462 => (x"e4",x"c0",x"51",x"66"),
  1463 => (x"81",x"c1",x"49",x"66"),
  1464 => (x"89",x"66",x"e0",x"c0"),
  1465 => (x"30",x"71",x"48",x"c1"),
  1466 => (x"89",x"c1",x"49",x"70"),
  1467 => (x"c3",x"7a",x"97",x"71"),
  1468 => (x"49",x"bf",x"ed",x"ca"),
  1469 => (x"29",x"66",x"e0",x"c0"),
  1470 => (x"48",x"4a",x"6a",x"97"),
  1471 => (x"f0",x"c0",x"98",x"71"),
  1472 => (x"49",x"6e",x"58",x"a6"),
  1473 => (x"4d",x"69",x"81",x"c4"),
  1474 => (x"d8",x"48",x"66",x"dc"),
  1475 => (x"c0",x"02",x"a8",x"66"),
  1476 => (x"a6",x"d8",x"87",x"c8"),
  1477 => (x"c0",x"78",x"c0",x"48"),
  1478 => (x"a6",x"d8",x"87",x"c5"),
  1479 => (x"d8",x"78",x"c1",x"48"),
  1480 => (x"e0",x"c0",x"1e",x"66"),
  1481 => (x"ff",x"49",x"75",x"1e"),
  1482 => (x"c8",x"87",x"e7",x"de"),
  1483 => (x"c0",x"4c",x"70",x"86"),
  1484 => (x"c1",x"06",x"ac",x"b7"),
  1485 => (x"85",x"74",x"87",x"d4"),
  1486 => (x"74",x"49",x"e0",x"c0"),
  1487 => (x"c1",x"4b",x"75",x"89"),
  1488 => (x"71",x"4a",x"c4",x"e1"),
  1489 => (x"87",x"e0",x"e5",x"fe"),
  1490 => (x"e8",x"c0",x"85",x"c2"),
  1491 => (x"80",x"c1",x"48",x"66"),
  1492 => (x"58",x"a6",x"ec",x"c0"),
  1493 => (x"49",x"66",x"ec",x"c0"),
  1494 => (x"a9",x"70",x"81",x"c1"),
  1495 => (x"87",x"c8",x"c0",x"02"),
  1496 => (x"c0",x"48",x"a6",x"d8"),
  1497 => (x"87",x"c5",x"c0",x"78"),
  1498 => (x"c1",x"48",x"a6",x"d8"),
  1499 => (x"1e",x"66",x"d8",x"78"),
  1500 => (x"c0",x"49",x"a4",x"c2"),
  1501 => (x"88",x"71",x"48",x"e0"),
  1502 => (x"75",x"1e",x"49",x"70"),
  1503 => (x"d1",x"dd",x"ff",x"49"),
  1504 => (x"c0",x"86",x"c8",x"87"),
  1505 => (x"ff",x"01",x"a8",x"b7"),
  1506 => (x"e8",x"c0",x"87",x"c0"),
  1507 => (x"d1",x"c0",x"02",x"66"),
  1508 => (x"c9",x"49",x"6e",x"87"),
  1509 => (x"66",x"e8",x"c0",x"81"),
  1510 => (x"c1",x"48",x"6e",x"51"),
  1511 => (x"c0",x"78",x"e6",x"cc"),
  1512 => (x"49",x"6e",x"87",x"cc"),
  1513 => (x"51",x"c2",x"81",x"c9"),
  1514 => (x"ef",x"c2",x"48",x"6e"),
  1515 => (x"7e",x"c1",x"78",x"e8"),
  1516 => (x"ff",x"87",x"c6",x"c0"),
  1517 => (x"70",x"87",x"c7",x"dc"),
  1518 => (x"c0",x"02",x"6e",x"4c"),
  1519 => (x"66",x"c4",x"87",x"f5"),
  1520 => (x"a8",x"66",x"c8",x"48"),
  1521 => (x"87",x"cb",x"c0",x"04"),
  1522 => (x"c1",x"48",x"66",x"c4"),
  1523 => (x"58",x"a6",x"c8",x"80"),
  1524 => (x"c8",x"87",x"e0",x"c0"),
  1525 => (x"88",x"c1",x"48",x"66"),
  1526 => (x"c0",x"58",x"a6",x"cc"),
  1527 => (x"c6",x"c1",x"87",x"d5"),
  1528 => (x"c8",x"c0",x"05",x"ac"),
  1529 => (x"48",x"66",x"cc",x"87"),
  1530 => (x"a6",x"d0",x"80",x"c1"),
  1531 => (x"cd",x"db",x"ff",x"58"),
  1532 => (x"d0",x"4c",x"70",x"87"),
  1533 => (x"80",x"c1",x"48",x"66"),
  1534 => (x"74",x"58",x"a6",x"d4"),
  1535 => (x"cb",x"c0",x"02",x"9c"),
  1536 => (x"48",x"66",x"c4",x"87"),
  1537 => (x"a8",x"66",x"c8",x"c1"),
  1538 => (x"87",x"ff",x"f2",x"04"),
  1539 => (x"87",x"e5",x"da",x"ff"),
  1540 => (x"c7",x"48",x"66",x"c4"),
  1541 => (x"e5",x"c0",x"03",x"a8"),
  1542 => (x"c0",x"c7",x"c3",x"87"),
  1543 => (x"c4",x"78",x"c0",x"48"),
  1544 => (x"91",x"cb",x"49",x"66"),
  1545 => (x"81",x"66",x"c0",x"c1"),
  1546 => (x"6a",x"4a",x"a1",x"c4"),
  1547 => (x"79",x"52",x"c0",x"4a"),
  1548 => (x"c1",x"48",x"66",x"c4"),
  1549 => (x"58",x"a6",x"c8",x"80"),
  1550 => (x"ff",x"04",x"a8",x"c7"),
  1551 => (x"d0",x"ff",x"87",x"db"),
  1552 => (x"87",x"cc",x"e1",x"8e"),
  1553 => (x"1e",x"00",x"20",x"3a"),
  1554 => (x"4b",x"71",x"1e",x"73"),
  1555 => (x"87",x"c6",x"02",x"9b"),
  1556 => (x"48",x"fc",x"c6",x"c3"),
  1557 => (x"1e",x"c7",x"78",x"c0"),
  1558 => (x"bf",x"fc",x"c6",x"c3"),
  1559 => (x"e4",x"c1",x"1e",x"49"),
  1560 => (x"c6",x"c3",x"1e",x"dc"),
  1561 => (x"ee",x"49",x"bf",x"f8"),
  1562 => (x"86",x"cc",x"87",x"f4"),
  1563 => (x"bf",x"f8",x"c6",x"c3"),
  1564 => (x"87",x"ca",x"ea",x"49"),
  1565 => (x"c8",x"02",x"9b",x"73"),
  1566 => (x"dc",x"e4",x"c1",x"87"),
  1567 => (x"f2",x"e5",x"c0",x"49"),
  1568 => (x"87",x"d0",x"e0",x"87"),
  1569 => (x"87",x"d6",x"c7",x"1e"),
  1570 => (x"fa",x"fe",x"49",x"c1"),
  1571 => (x"cf",x"ea",x"fe",x"87"),
  1572 => (x"02",x"98",x"70",x"87"),
  1573 => (x"f3",x"fe",x"87",x"cd"),
  1574 => (x"98",x"70",x"87",x"cc"),
  1575 => (x"c1",x"87",x"c4",x"02"),
  1576 => (x"c0",x"87",x"c2",x"4a"),
  1577 => (x"05",x"9a",x"72",x"4a"),
  1578 => (x"1e",x"c0",x"87",x"ce"),
  1579 => (x"49",x"d5",x"e3",x"c1"),
  1580 => (x"87",x"c4",x"f1",x"c0"),
  1581 => (x"87",x"fe",x"86",x"c4"),
  1582 => (x"e3",x"c1",x"1e",x"c0"),
  1583 => (x"f0",x"c0",x"49",x"e0"),
  1584 => (x"1e",x"c0",x"87",x"f6"),
  1585 => (x"87",x"e7",x"d1",x"c1"),
  1586 => (x"f0",x"c0",x"49",x"70"),
  1587 => (x"cc",x"c3",x"87",x"ea"),
  1588 => (x"26",x"8e",x"f8",x"87"),
  1589 => (x"20",x"44",x"53",x"4f"),
  1590 => (x"6c",x"69",x"61",x"66"),
  1591 => (x"00",x"2e",x"64",x"65"),
  1592 => (x"74",x"6f",x"6f",x"42"),
  1593 => (x"2e",x"67",x"6e",x"69"),
  1594 => (x"1e",x"00",x"2e",x"2e"),
  1595 => (x"87",x"d2",x"e8",x"c0"),
  1596 => (x"87",x"fa",x"f3",x"c0"),
  1597 => (x"4f",x"26",x"87",x"f6"),
  1598 => (x"fc",x"c6",x"c3",x"1e"),
  1599 => (x"c3",x"78",x"c0",x"48"),
  1600 => (x"c0",x"48",x"f8",x"c6"),
  1601 => (x"87",x"fc",x"fd",x"78"),
  1602 => (x"48",x"c0",x"87",x"e1"),
  1603 => (x"20",x"80",x"4f",x"26"),
  1604 => (x"74",x"69",x"78",x"45"),
  1605 => (x"42",x"20",x"80",x"00"),
  1606 => (x"00",x"6b",x"63",x"61"),
  1607 => (x"00",x"00",x"12",x"d6"),
  1608 => (x"00",x"00",x"31",x"d1"),
  1609 => (x"d6",x"00",x"00",x"00"),
  1610 => (x"ef",x"00",x"00",x"12"),
  1611 => (x"00",x"00",x"00",x"31"),
  1612 => (x"12",x"d6",x"00",x"00"),
  1613 => (x"32",x"0d",x"00",x"00"),
  1614 => (x"00",x"00",x"00",x"00"),
  1615 => (x"00",x"12",x"d6",x"00"),
  1616 => (x"00",x"32",x"2b",x"00"),
  1617 => (x"00",x"00",x"00",x"00"),
  1618 => (x"00",x"00",x"12",x"d6"),
  1619 => (x"00",x"00",x"32",x"49"),
  1620 => (x"d6",x"00",x"00",x"00"),
  1621 => (x"67",x"00",x"00",x"12"),
  1622 => (x"00",x"00",x"00",x"32"),
  1623 => (x"12",x"d6",x"00",x"00"),
  1624 => (x"32",x"85",x"00",x"00"),
  1625 => (x"00",x"00",x"00",x"00"),
  1626 => (x"00",x"12",x"d6",x"00"),
  1627 => (x"00",x"00",x"00",x"00"),
  1628 => (x"00",x"00",x"00",x"00"),
  1629 => (x"00",x"00",x"13",x"5a"),
  1630 => (x"00",x"00",x"00",x"00"),
  1631 => (x"4c",x"00",x"00",x"00"),
  1632 => (x"20",x"64",x"61",x"6f"),
  1633 => (x"1e",x"00",x"2e",x"2a"),
  1634 => (x"c0",x"48",x"f0",x"fe"),
  1635 => (x"79",x"09",x"cd",x"78"),
  1636 => (x"1e",x"4f",x"26",x"09"),
  1637 => (x"bf",x"f0",x"fe",x"1e"),
  1638 => (x"26",x"26",x"48",x"7e"),
  1639 => (x"f0",x"fe",x"1e",x"4f"),
  1640 => (x"26",x"78",x"c1",x"48"),
  1641 => (x"f0",x"fe",x"1e",x"4f"),
  1642 => (x"26",x"78",x"c0",x"48"),
  1643 => (x"4a",x"71",x"1e",x"4f"),
  1644 => (x"26",x"52",x"52",x"c0"),
  1645 => (x"5b",x"5e",x"0e",x"4f"),
  1646 => (x"f4",x"0e",x"5d",x"5c"),
  1647 => (x"97",x"4d",x"71",x"86"),
  1648 => (x"a5",x"c1",x"7e",x"6d"),
  1649 => (x"48",x"6c",x"97",x"4c"),
  1650 => (x"6e",x"58",x"a6",x"c8"),
  1651 => (x"a8",x"66",x"c4",x"48"),
  1652 => (x"ff",x"87",x"c5",x"05"),
  1653 => (x"87",x"e6",x"c0",x"48"),
  1654 => (x"c2",x"87",x"ca",x"ff"),
  1655 => (x"6c",x"97",x"49",x"a5"),
  1656 => (x"4b",x"a3",x"71",x"4b"),
  1657 => (x"97",x"4b",x"6b",x"97"),
  1658 => (x"48",x"6e",x"7e",x"6c"),
  1659 => (x"a6",x"c8",x"80",x"c1"),
  1660 => (x"cc",x"98",x"c7",x"58"),
  1661 => (x"97",x"70",x"58",x"a6"),
  1662 => (x"87",x"e1",x"fe",x"7c"),
  1663 => (x"8e",x"f4",x"48",x"73"),
  1664 => (x"4c",x"26",x"4d",x"26"),
  1665 => (x"4f",x"26",x"4b",x"26"),
  1666 => (x"5c",x"5b",x"5e",x"0e"),
  1667 => (x"71",x"86",x"f4",x"0e"),
  1668 => (x"4a",x"66",x"d8",x"4c"),
  1669 => (x"c2",x"9a",x"ff",x"c3"),
  1670 => (x"6c",x"97",x"4b",x"a4"),
  1671 => (x"49",x"a1",x"73",x"49"),
  1672 => (x"6c",x"97",x"51",x"72"),
  1673 => (x"c1",x"48",x"6e",x"7e"),
  1674 => (x"58",x"a6",x"c8",x"80"),
  1675 => (x"a6",x"cc",x"98",x"c7"),
  1676 => (x"f4",x"54",x"70",x"58"),
  1677 => (x"87",x"ca",x"ff",x"8e"),
  1678 => (x"e8",x"fd",x"1e",x"1e"),
  1679 => (x"4a",x"bf",x"e0",x"87"),
  1680 => (x"c0",x"e0",x"c0",x"49"),
  1681 => (x"87",x"cb",x"02",x"99"),
  1682 => (x"ca",x"c3",x"1e",x"72"),
  1683 => (x"f7",x"fe",x"49",x"e3"),
  1684 => (x"fc",x"86",x"c4",x"87"),
  1685 => (x"7e",x"70",x"87",x"fd"),
  1686 => (x"26",x"87",x"c2",x"fd"),
  1687 => (x"c3",x"1e",x"4f",x"26"),
  1688 => (x"fd",x"49",x"e3",x"ca"),
  1689 => (x"e8",x"c1",x"87",x"c7"),
  1690 => (x"da",x"fc",x"49",x"f8"),
  1691 => (x"87",x"d0",x"c5",x"87"),
  1692 => (x"5e",x"0e",x"4f",x"26"),
  1693 => (x"0e",x"5d",x"5c",x"5b"),
  1694 => (x"bf",x"c2",x"cb",x"c3"),
  1695 => (x"c6",x"eb",x"c1",x"4a"),
  1696 => (x"72",x"4c",x"49",x"bf"),
  1697 => (x"fc",x"4d",x"71",x"bc"),
  1698 => (x"4b",x"c0",x"87",x"db"),
  1699 => (x"99",x"d0",x"49",x"74"),
  1700 => (x"75",x"87",x"d5",x"02"),
  1701 => (x"71",x"99",x"d0",x"49"),
  1702 => (x"c1",x"1e",x"c0",x"1e"),
  1703 => (x"73",x"4a",x"cf",x"f1"),
  1704 => (x"c0",x"49",x"12",x"82"),
  1705 => (x"86",x"c8",x"87",x"e4"),
  1706 => (x"83",x"2d",x"2c",x"c1"),
  1707 => (x"ff",x"04",x"ab",x"c8"),
  1708 => (x"e8",x"fb",x"87",x"da"),
  1709 => (x"c6",x"eb",x"c1",x"87"),
  1710 => (x"c2",x"cb",x"c3",x"48"),
  1711 => (x"4d",x"26",x"78",x"bf"),
  1712 => (x"4b",x"26",x"4c",x"26"),
  1713 => (x"00",x"00",x"4f",x"26"),
  1714 => (x"ff",x"1e",x"00",x"00"),
  1715 => (x"e1",x"c8",x"48",x"d0"),
  1716 => (x"48",x"d4",x"ff",x"78"),
  1717 => (x"66",x"c4",x"78",x"c5"),
  1718 => (x"c3",x"87",x"c3",x"02"),
  1719 => (x"66",x"c8",x"78",x"e0"),
  1720 => (x"ff",x"87",x"c6",x"02"),
  1721 => (x"f0",x"c3",x"48",x"d4"),
  1722 => (x"48",x"d4",x"ff",x"78"),
  1723 => (x"d0",x"ff",x"78",x"71"),
  1724 => (x"78",x"e1",x"c8",x"48"),
  1725 => (x"26",x"78",x"e0",x"c0"),
  1726 => (x"5b",x"5e",x"0e",x"4f"),
  1727 => (x"4c",x"71",x"0e",x"5c"),
  1728 => (x"49",x"e3",x"ca",x"c3"),
  1729 => (x"70",x"87",x"ee",x"fa"),
  1730 => (x"aa",x"b7",x"c0",x"4a"),
  1731 => (x"87",x"e3",x"c2",x"04"),
  1732 => (x"05",x"aa",x"e0",x"c3"),
  1733 => (x"ee",x"c1",x"87",x"c9"),
  1734 => (x"78",x"c1",x"48",x"fc"),
  1735 => (x"c3",x"87",x"d4",x"c2"),
  1736 => (x"c9",x"05",x"aa",x"f0"),
  1737 => (x"f8",x"ee",x"c1",x"87"),
  1738 => (x"c1",x"78",x"c1",x"48"),
  1739 => (x"ee",x"c1",x"87",x"f5"),
  1740 => (x"c7",x"02",x"bf",x"fc"),
  1741 => (x"c2",x"4b",x"72",x"87"),
  1742 => (x"87",x"c2",x"b3",x"c0"),
  1743 => (x"9c",x"74",x"4b",x"72"),
  1744 => (x"c1",x"87",x"d1",x"05"),
  1745 => (x"1e",x"bf",x"f8",x"ee"),
  1746 => (x"bf",x"fc",x"ee",x"c1"),
  1747 => (x"fd",x"49",x"72",x"1e"),
  1748 => (x"86",x"c8",x"87",x"f8"),
  1749 => (x"bf",x"f8",x"ee",x"c1"),
  1750 => (x"87",x"e0",x"c0",x"02"),
  1751 => (x"b7",x"c4",x"49",x"73"),
  1752 => (x"f0",x"c1",x"91",x"29"),
  1753 => (x"4a",x"73",x"81",x"cf"),
  1754 => (x"92",x"c2",x"9a",x"cf"),
  1755 => (x"30",x"72",x"48",x"c1"),
  1756 => (x"ba",x"ff",x"4a",x"70"),
  1757 => (x"98",x"69",x"48",x"72"),
  1758 => (x"87",x"db",x"79",x"70"),
  1759 => (x"b7",x"c4",x"49",x"73"),
  1760 => (x"f0",x"c1",x"91",x"29"),
  1761 => (x"4a",x"73",x"81",x"cf"),
  1762 => (x"92",x"c2",x"9a",x"cf"),
  1763 => (x"30",x"72",x"48",x"c3"),
  1764 => (x"69",x"48",x"4a",x"70"),
  1765 => (x"c1",x"79",x"70",x"b0"),
  1766 => (x"c0",x"48",x"fc",x"ee"),
  1767 => (x"f8",x"ee",x"c1",x"78"),
  1768 => (x"c3",x"78",x"c0",x"48"),
  1769 => (x"f8",x"49",x"e3",x"ca"),
  1770 => (x"4a",x"70",x"87",x"cb"),
  1771 => (x"03",x"aa",x"b7",x"c0"),
  1772 => (x"c0",x"87",x"dd",x"fd"),
  1773 => (x"87",x"c8",x"fc",x"48"),
  1774 => (x"00",x"00",x"00",x"00"),
  1775 => (x"00",x"00",x"00",x"00"),
  1776 => (x"72",x"4a",x"c0",x"1e"),
  1777 => (x"c1",x"91",x"c4",x"49"),
  1778 => (x"c0",x"81",x"cf",x"f0"),
  1779 => (x"d0",x"82",x"c1",x"79"),
  1780 => (x"ee",x"04",x"aa",x"b7"),
  1781 => (x"0e",x"4f",x"26",x"87"),
  1782 => (x"5d",x"5c",x"5b",x"5e"),
  1783 => (x"f7",x"4d",x"71",x"0e"),
  1784 => (x"4a",x"75",x"87",x"c3"),
  1785 => (x"92",x"2a",x"b7",x"c4"),
  1786 => (x"82",x"cf",x"f0",x"c1"),
  1787 => (x"9c",x"cf",x"4c",x"75"),
  1788 => (x"49",x"6a",x"94",x"c2"),
  1789 => (x"c3",x"2b",x"74",x"4b"),
  1790 => (x"74",x"48",x"c2",x"9b"),
  1791 => (x"ff",x"4c",x"70",x"30"),
  1792 => (x"71",x"48",x"74",x"bc"),
  1793 => (x"f6",x"7a",x"70",x"98"),
  1794 => (x"48",x"73",x"87",x"d3"),
  1795 => (x"00",x"87",x"ef",x"fa"),
  1796 => (x"00",x"00",x"00",x"00"),
  1797 => (x"00",x"00",x"00",x"00"),
  1798 => (x"00",x"00",x"00",x"00"),
  1799 => (x"00",x"00",x"00",x"00"),
  1800 => (x"00",x"00",x"00",x"00"),
  1801 => (x"00",x"00",x"00",x"00"),
  1802 => (x"00",x"00",x"00",x"00"),
  1803 => (x"00",x"00",x"00",x"00"),
  1804 => (x"00",x"00",x"00",x"00"),
  1805 => (x"00",x"00",x"00",x"00"),
  1806 => (x"00",x"00",x"00",x"00"),
  1807 => (x"00",x"00",x"00",x"00"),
  1808 => (x"00",x"00",x"00",x"00"),
  1809 => (x"00",x"00",x"00",x"00"),
  1810 => (x"00",x"00",x"00",x"00"),
  1811 => (x"16",x"00",x"00",x"00"),
  1812 => (x"2e",x"25",x"26",x"1e"),
  1813 => (x"1e",x"3e",x"3d",x"36"),
  1814 => (x"c8",x"48",x"d0",x"ff"),
  1815 => (x"48",x"71",x"78",x"e1"),
  1816 => (x"78",x"08",x"d4",x"ff"),
  1817 => (x"ff",x"1e",x"4f",x"26"),
  1818 => (x"e1",x"c8",x"48",x"d0"),
  1819 => (x"ff",x"48",x"71",x"78"),
  1820 => (x"c4",x"78",x"08",x"d4"),
  1821 => (x"d4",x"ff",x"48",x"66"),
  1822 => (x"4f",x"26",x"78",x"08"),
  1823 => (x"c4",x"4a",x"71",x"1e"),
  1824 => (x"72",x"1e",x"49",x"66"),
  1825 => (x"87",x"de",x"ff",x"49"),
  1826 => (x"c0",x"48",x"d0",x"ff"),
  1827 => (x"26",x"26",x"78",x"e0"),
  1828 => (x"4a",x"71",x"1e",x"4f"),
  1829 => (x"c1",x"1e",x"66",x"c4"),
  1830 => (x"ff",x"49",x"a2",x"e0"),
  1831 => (x"66",x"c8",x"87",x"c8"),
  1832 => (x"29",x"b7",x"c8",x"49"),
  1833 => (x"71",x"48",x"d4",x"ff"),
  1834 => (x"48",x"d0",x"ff",x"78"),
  1835 => (x"26",x"78",x"e0",x"c0"),
  1836 => (x"71",x"1e",x"4f",x"26"),
  1837 => (x"49",x"da",x"1e",x"4a"),
  1838 => (x"c8",x"87",x"eb",x"fe"),
  1839 => (x"c8",x"49",x"bf",x"66"),
  1840 => (x"80",x"c4",x"48",x"66"),
  1841 => (x"c8",x"58",x"a6",x"cc"),
  1842 => (x"d4",x"ff",x"29",x"b7"),
  1843 => (x"c8",x"78",x"71",x"48"),
  1844 => (x"c8",x"49",x"bf",x"66"),
  1845 => (x"78",x"71",x"29",x"b7"),
  1846 => (x"c0",x"48",x"d0",x"ff"),
  1847 => (x"26",x"26",x"78",x"e0"),
  1848 => (x"d4",x"ff",x"1e",x"4f"),
  1849 => (x"7a",x"ff",x"c3",x"4a"),
  1850 => (x"c8",x"48",x"d0",x"ff"),
  1851 => (x"7a",x"de",x"78",x"e1"),
  1852 => (x"bf",x"ed",x"ca",x"c3"),
  1853 => (x"c8",x"48",x"49",x"7a"),
  1854 => (x"71",x"7a",x"70",x"28"),
  1855 => (x"70",x"28",x"d0",x"48"),
  1856 => (x"d8",x"48",x"71",x"7a"),
  1857 => (x"ff",x"7a",x"70",x"28"),
  1858 => (x"e0",x"c0",x"48",x"d0"),
  1859 => (x"0e",x"4f",x"26",x"78"),
  1860 => (x"5d",x"5c",x"5b",x"5e"),
  1861 => (x"c3",x"4c",x"71",x"0e"),
  1862 => (x"4d",x"bf",x"ed",x"ca"),
  1863 => (x"d0",x"2b",x"74",x"4b"),
  1864 => (x"83",x"c1",x"9b",x"66"),
  1865 => (x"04",x"ab",x"66",x"d4"),
  1866 => (x"4b",x"c0",x"87",x"c2"),
  1867 => (x"66",x"d0",x"4a",x"74"),
  1868 => (x"ff",x"31",x"72",x"49"),
  1869 => (x"73",x"99",x"75",x"b9"),
  1870 => (x"70",x"30",x"72",x"48"),
  1871 => (x"b0",x"71",x"48",x"4a"),
  1872 => (x"58",x"f1",x"ca",x"c3"),
  1873 => (x"26",x"87",x"da",x"fe"),
  1874 => (x"26",x"4c",x"26",x"4d"),
  1875 => (x"1e",x"4f",x"26",x"4b"),
  1876 => (x"c8",x"48",x"d0",x"ff"),
  1877 => (x"48",x"71",x"78",x"c9"),
  1878 => (x"78",x"08",x"d4",x"ff"),
  1879 => (x"71",x"1e",x"4f",x"26"),
  1880 => (x"87",x"eb",x"49",x"4a"),
  1881 => (x"c8",x"48",x"d0",x"ff"),
  1882 => (x"1e",x"4f",x"26",x"78"),
  1883 => (x"4b",x"71",x"1e",x"73"),
  1884 => (x"bf",x"fd",x"ca",x"c3"),
  1885 => (x"c2",x"87",x"c3",x"02"),
  1886 => (x"d0",x"ff",x"87",x"eb"),
  1887 => (x"78",x"c9",x"c8",x"48"),
  1888 => (x"e0",x"c0",x"49",x"73"),
  1889 => (x"48",x"d4",x"ff",x"b1"),
  1890 => (x"ca",x"c3",x"78",x"71"),
  1891 => (x"78",x"c0",x"48",x"f1"),
  1892 => (x"c5",x"02",x"66",x"c8"),
  1893 => (x"49",x"ff",x"c3",x"87"),
  1894 => (x"49",x"c0",x"87",x"c2"),
  1895 => (x"59",x"f9",x"ca",x"c3"),
  1896 => (x"c6",x"02",x"66",x"cc"),
  1897 => (x"d5",x"d5",x"c5",x"87"),
  1898 => (x"cf",x"87",x"c4",x"4a"),
  1899 => (x"c3",x"4a",x"ff",x"ff"),
  1900 => (x"c3",x"5a",x"fd",x"ca"),
  1901 => (x"c1",x"48",x"fd",x"ca"),
  1902 => (x"26",x"87",x"c4",x"78"),
  1903 => (x"26",x"4c",x"26",x"4d"),
  1904 => (x"0e",x"4f",x"26",x"4b"),
  1905 => (x"5d",x"5c",x"5b",x"5e"),
  1906 => (x"c3",x"4a",x"71",x"0e"),
  1907 => (x"4c",x"bf",x"f9",x"ca"),
  1908 => (x"cb",x"02",x"9a",x"72"),
  1909 => (x"91",x"c8",x"49",x"87"),
  1910 => (x"4b",x"e1",x"f5",x"c1"),
  1911 => (x"87",x"c4",x"83",x"71"),
  1912 => (x"4b",x"e1",x"f9",x"c1"),
  1913 => (x"49",x"13",x"4d",x"c0"),
  1914 => (x"ca",x"c3",x"99",x"74"),
  1915 => (x"ff",x"b9",x"bf",x"f5"),
  1916 => (x"78",x"71",x"48",x"d4"),
  1917 => (x"85",x"2c",x"b7",x"c1"),
  1918 => (x"04",x"ad",x"b7",x"c8"),
  1919 => (x"ca",x"c3",x"87",x"e8"),
  1920 => (x"c8",x"48",x"bf",x"f1"),
  1921 => (x"f5",x"ca",x"c3",x"80"),
  1922 => (x"87",x"ef",x"fe",x"58"),
  1923 => (x"71",x"1e",x"73",x"1e"),
  1924 => (x"9a",x"4a",x"13",x"4b"),
  1925 => (x"72",x"87",x"cb",x"02"),
  1926 => (x"87",x"e7",x"fe",x"49"),
  1927 => (x"05",x"9a",x"4a",x"13"),
  1928 => (x"da",x"fe",x"87",x"f5"),
  1929 => (x"ca",x"c3",x"1e",x"87"),
  1930 => (x"c3",x"49",x"bf",x"f1"),
  1931 => (x"c1",x"48",x"f1",x"ca"),
  1932 => (x"c0",x"c4",x"78",x"a1"),
  1933 => (x"db",x"03",x"a9",x"b7"),
  1934 => (x"48",x"d4",x"ff",x"87"),
  1935 => (x"bf",x"f5",x"ca",x"c3"),
  1936 => (x"f1",x"ca",x"c3",x"78"),
  1937 => (x"ca",x"c3",x"49",x"bf"),
  1938 => (x"a1",x"c1",x"48",x"f1"),
  1939 => (x"b7",x"c0",x"c4",x"78"),
  1940 => (x"87",x"e5",x"04",x"a9"),
  1941 => (x"c8",x"48",x"d0",x"ff"),
  1942 => (x"fd",x"ca",x"c3",x"78"),
  1943 => (x"26",x"78",x"c0",x"48"),
  1944 => (x"00",x"00",x"00",x"4f"),
  1945 => (x"00",x"00",x"00",x"00"),
  1946 => (x"00",x"00",x"00",x"00"),
  1947 => (x"00",x"00",x"5f",x"5f"),
  1948 => (x"03",x"03",x"00",x"00"),
  1949 => (x"00",x"03",x"03",x"00"),
  1950 => (x"7f",x"7f",x"14",x"00"),
  1951 => (x"14",x"7f",x"7f",x"14"),
  1952 => (x"2e",x"24",x"00",x"00"),
  1953 => (x"12",x"3a",x"6b",x"6b"),
  1954 => (x"36",x"6a",x"4c",x"00"),
  1955 => (x"32",x"56",x"6c",x"18"),
  1956 => (x"4f",x"7e",x"30",x"00"),
  1957 => (x"68",x"3a",x"77",x"59"),
  1958 => (x"04",x"00",x"00",x"40"),
  1959 => (x"00",x"00",x"03",x"07"),
  1960 => (x"1c",x"00",x"00",x"00"),
  1961 => (x"00",x"41",x"63",x"3e"),
  1962 => (x"41",x"00",x"00",x"00"),
  1963 => (x"00",x"1c",x"3e",x"63"),
  1964 => (x"3e",x"2a",x"08",x"00"),
  1965 => (x"2a",x"3e",x"1c",x"1c"),
  1966 => (x"08",x"08",x"00",x"08"),
  1967 => (x"08",x"08",x"3e",x"3e"),
  1968 => (x"80",x"00",x"00",x"00"),
  1969 => (x"00",x"00",x"60",x"e0"),
  1970 => (x"08",x"08",x"00",x"00"),
  1971 => (x"08",x"08",x"08",x"08"),
  1972 => (x"00",x"00",x"00",x"00"),
  1973 => (x"00",x"00",x"60",x"60"),
  1974 => (x"30",x"60",x"40",x"00"),
  1975 => (x"03",x"06",x"0c",x"18"),
  1976 => (x"7f",x"3e",x"00",x"01"),
  1977 => (x"3e",x"7f",x"4d",x"59"),
  1978 => (x"06",x"04",x"00",x"00"),
  1979 => (x"00",x"00",x"7f",x"7f"),
  1980 => (x"63",x"42",x"00",x"00"),
  1981 => (x"46",x"4f",x"59",x"71"),
  1982 => (x"63",x"22",x"00",x"00"),
  1983 => (x"36",x"7f",x"49",x"49"),
  1984 => (x"16",x"1c",x"18",x"00"),
  1985 => (x"10",x"7f",x"7f",x"13"),
  1986 => (x"67",x"27",x"00",x"00"),
  1987 => (x"39",x"7d",x"45",x"45"),
  1988 => (x"7e",x"3c",x"00",x"00"),
  1989 => (x"30",x"79",x"49",x"4b"),
  1990 => (x"01",x"01",x"00",x"00"),
  1991 => (x"07",x"0f",x"79",x"71"),
  1992 => (x"7f",x"36",x"00",x"00"),
  1993 => (x"36",x"7f",x"49",x"49"),
  1994 => (x"4f",x"06",x"00",x"00"),
  1995 => (x"1e",x"3f",x"69",x"49"),
  1996 => (x"00",x"00",x"00",x"00"),
  1997 => (x"00",x"00",x"66",x"66"),
  1998 => (x"80",x"00",x"00",x"00"),
  1999 => (x"00",x"00",x"66",x"e6"),
  2000 => (x"08",x"08",x"00",x"00"),
  2001 => (x"22",x"22",x"14",x"14"),
  2002 => (x"14",x"14",x"00",x"00"),
  2003 => (x"14",x"14",x"14",x"14"),
  2004 => (x"22",x"22",x"00",x"00"),
  2005 => (x"08",x"08",x"14",x"14"),
  2006 => (x"03",x"02",x"00",x"00"),
  2007 => (x"06",x"0f",x"59",x"51"),
  2008 => (x"41",x"7f",x"3e",x"00"),
  2009 => (x"1e",x"1f",x"55",x"5d"),
  2010 => (x"7f",x"7e",x"00",x"00"),
  2011 => (x"7e",x"7f",x"09",x"09"),
  2012 => (x"7f",x"7f",x"00",x"00"),
  2013 => (x"36",x"7f",x"49",x"49"),
  2014 => (x"3e",x"1c",x"00",x"00"),
  2015 => (x"41",x"41",x"41",x"63"),
  2016 => (x"7f",x"7f",x"00",x"00"),
  2017 => (x"1c",x"3e",x"63",x"41"),
  2018 => (x"7f",x"7f",x"00",x"00"),
  2019 => (x"41",x"41",x"49",x"49"),
  2020 => (x"7f",x"7f",x"00",x"00"),
  2021 => (x"01",x"01",x"09",x"09"),
  2022 => (x"7f",x"3e",x"00",x"00"),
  2023 => (x"7a",x"7b",x"49",x"41"),
  2024 => (x"7f",x"7f",x"00",x"00"),
  2025 => (x"7f",x"7f",x"08",x"08"),
  2026 => (x"41",x"00",x"00",x"00"),
  2027 => (x"00",x"41",x"7f",x"7f"),
  2028 => (x"60",x"20",x"00",x"00"),
  2029 => (x"3f",x"7f",x"40",x"40"),
  2030 => (x"08",x"7f",x"7f",x"00"),
  2031 => (x"41",x"63",x"36",x"1c"),
  2032 => (x"7f",x"7f",x"00",x"00"),
  2033 => (x"40",x"40",x"40",x"40"),
  2034 => (x"06",x"7f",x"7f",x"00"),
  2035 => (x"7f",x"7f",x"06",x"0c"),
  2036 => (x"06",x"7f",x"7f",x"00"),
  2037 => (x"7f",x"7f",x"18",x"0c"),
  2038 => (x"7f",x"3e",x"00",x"00"),
  2039 => (x"3e",x"7f",x"41",x"41"),
  2040 => (x"7f",x"7f",x"00",x"00"),
  2041 => (x"06",x"0f",x"09",x"09"),
  2042 => (x"41",x"7f",x"3e",x"00"),
  2043 => (x"40",x"7e",x"7f",x"61"),
  2044 => (x"7f",x"7f",x"00",x"00"),
  2045 => (x"66",x"7f",x"19",x"09"),
  2046 => (x"6f",x"26",x"00",x"00"),
  2047 => (x"32",x"7b",x"59",x"4d"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

