`define DEMISTIFY
`define VIVADO
