
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"4b",x"26",x"4c",x"26"),
     1 => (x"71",x"1e",x"4f",x"26"),
     2 => (x"d2",x"ee",x"c2",x"4a"),
     3 => (x"d2",x"ee",x"c2",x"5a"),
     4 => (x"49",x"78",x"c7",x"48"),
     5 => (x"26",x"87",x"dd",x"fe"),
     6 => (x"1e",x"73",x"1e",x"4f"),
     7 => (x"b7",x"c0",x"4a",x"71"),
     8 => (x"87",x"d3",x"03",x"aa"),
     9 => (x"bf",x"f0",x"ce",x"c2"),
    10 => (x"c1",x"87",x"c4",x"05"),
    11 => (x"c0",x"87",x"c2",x"4b"),
    12 => (x"f4",x"ce",x"c2",x"4b"),
    13 => (x"c2",x"87",x"c4",x"5b"),
    14 => (x"c2",x"5a",x"f4",x"ce"),
    15 => (x"4a",x"bf",x"f0",x"ce"),
    16 => (x"c0",x"c1",x"9a",x"c1"),
    17 => (x"e8",x"ec",x"49",x"a2"),
    18 => (x"c2",x"48",x"fc",x"87"),
    19 => (x"78",x"bf",x"f0",x"ce"),
    20 => (x"1e",x"87",x"ef",x"fe"),
    21 => (x"66",x"c4",x"4a",x"71"),
    22 => (x"e9",x"49",x"72",x"1e"),
    23 => (x"26",x"26",x"87",x"f5"),
    24 => (x"ce",x"c2",x"1e",x"4f"),
    25 => (x"e6",x"49",x"bf",x"f0"),
    26 => (x"ee",x"c2",x"87",x"cf"),
    27 => (x"bf",x"e8",x"48",x"c6"),
    28 => (x"c2",x"ee",x"c2",x"78"),
    29 => (x"78",x"bf",x"ec",x"48"),
    30 => (x"bf",x"c6",x"ee",x"c2"),
    31 => (x"ff",x"c3",x"49",x"4a"),
    32 => (x"2a",x"b7",x"c8",x"99"),
    33 => (x"b0",x"71",x"48",x"72"),
    34 => (x"58",x"ce",x"ee",x"c2"),
    35 => (x"5e",x"0e",x"4f",x"26"),
    36 => (x"0e",x"5d",x"5c",x"5b"),
    37 => (x"c8",x"ff",x"4b",x"71"),
    38 => (x"c1",x"ee",x"c2",x"87"),
    39 => (x"73",x"50",x"c0",x"48"),
    40 => (x"87",x"f5",x"e5",x"49"),
    41 => (x"c2",x"4c",x"49",x"70"),
    42 => (x"49",x"ee",x"cb",x"9c"),
    43 => (x"70",x"87",x"c9",x"cc"),
    44 => (x"ee",x"c2",x"4d",x"49"),
    45 => (x"05",x"bf",x"97",x"c1"),
    46 => (x"d0",x"87",x"e2",x"c1"),
    47 => (x"ee",x"c2",x"49",x"66"),
    48 => (x"05",x"99",x"bf",x"ca"),
    49 => (x"66",x"d4",x"87",x"d6"),
    50 => (x"c2",x"ee",x"c2",x"49"),
    51 => (x"cb",x"05",x"99",x"bf"),
    52 => (x"e5",x"49",x"73",x"87"),
    53 => (x"98",x"70",x"87",x"c3"),
    54 => (x"87",x"c1",x"c1",x"02"),
    55 => (x"c0",x"fe",x"4c",x"c1"),
    56 => (x"cb",x"49",x"75",x"87"),
    57 => (x"98",x"70",x"87",x"de"),
    58 => (x"c2",x"87",x"c6",x"02"),
    59 => (x"c1",x"48",x"c1",x"ee"),
    60 => (x"c1",x"ee",x"c2",x"50"),
    61 => (x"c0",x"05",x"bf",x"97"),
    62 => (x"ee",x"c2",x"87",x"e3"),
    63 => (x"d0",x"49",x"bf",x"ca"),
    64 => (x"ff",x"05",x"99",x"66"),
    65 => (x"ee",x"c2",x"87",x"d6"),
    66 => (x"d4",x"49",x"bf",x"c2"),
    67 => (x"ff",x"05",x"99",x"66"),
    68 => (x"49",x"73",x"87",x"ca"),
    69 => (x"70",x"87",x"c2",x"e4"),
    70 => (x"ff",x"fe",x"05",x"98"),
    71 => (x"fb",x"48",x"74",x"87"),
    72 => (x"5e",x"0e",x"87",x"dc"),
    73 => (x"0e",x"5d",x"5c",x"5b"),
    74 => (x"4d",x"c0",x"86",x"f4"),
    75 => (x"7e",x"bf",x"ec",x"4c"),
    76 => (x"c2",x"48",x"a6",x"c4"),
    77 => (x"78",x"bf",x"ce",x"ee"),
    78 => (x"1e",x"c0",x"1e",x"c1"),
    79 => (x"cd",x"fd",x"49",x"c7"),
    80 => (x"70",x"86",x"c8",x"87"),
    81 => (x"87",x"cd",x"02",x"98"),
    82 => (x"cc",x"fb",x"49",x"ff"),
    83 => (x"49",x"da",x"c1",x"87"),
    84 => (x"c1",x"87",x"c6",x"e3"),
    85 => (x"c1",x"ee",x"c2",x"4d"),
    86 => (x"c3",x"02",x"bf",x"97"),
    87 => (x"87",x"ee",x"d5",x"87"),
    88 => (x"bf",x"c6",x"ee",x"c2"),
    89 => (x"f0",x"ce",x"c2",x"4b"),
    90 => (x"d9",x"c1",x"05",x"bf"),
    91 => (x"48",x"a6",x"c4",x"87"),
    92 => (x"78",x"c0",x"c0",x"c8"),
    93 => (x"7e",x"dc",x"ce",x"c2"),
    94 => (x"49",x"bf",x"97",x"6e"),
    95 => (x"80",x"c1",x"48",x"6e"),
    96 => (x"e2",x"71",x"7e",x"70"),
    97 => (x"98",x"70",x"87",x"d3"),
    98 => (x"c4",x"87",x"c3",x"02"),
    99 => (x"66",x"c4",x"b3",x"66"),
   100 => (x"28",x"b7",x"c1",x"48"),
   101 => (x"70",x"58",x"a6",x"c8"),
   102 => (x"db",x"ff",x"05",x"98"),
   103 => (x"49",x"fd",x"c3",x"87"),
   104 => (x"c3",x"87",x"f6",x"e1"),
   105 => (x"f0",x"e1",x"49",x"fa"),
   106 => (x"c3",x"49",x"73",x"87"),
   107 => (x"1e",x"71",x"99",x"ff"),
   108 => (x"de",x"fa",x"49",x"c0"),
   109 => (x"c8",x"49",x"73",x"87"),
   110 => (x"1e",x"71",x"29",x"b7"),
   111 => (x"d2",x"fa",x"49",x"c1"),
   112 => (x"c5",x"86",x"c8",x"87"),
   113 => (x"ee",x"c2",x"87",x"ff"),
   114 => (x"9b",x"4b",x"bf",x"ca"),
   115 => (x"c2",x"87",x"dd",x"02"),
   116 => (x"49",x"bf",x"ec",x"ce"),
   117 => (x"70",x"87",x"ed",x"c7"),
   118 => (x"87",x"c4",x"05",x"98"),
   119 => (x"87",x"d2",x"4b",x"c0"),
   120 => (x"c7",x"49",x"e0",x"c2"),
   121 => (x"ce",x"c2",x"87",x"d2"),
   122 => (x"87",x"c6",x"58",x"f0"),
   123 => (x"48",x"ec",x"ce",x"c2"),
   124 => (x"49",x"73",x"78",x"c0"),
   125 => (x"cd",x"05",x"99",x"c2"),
   126 => (x"49",x"eb",x"c3",x"87"),
   127 => (x"70",x"87",x"da",x"e0"),
   128 => (x"02",x"99",x"c2",x"49"),
   129 => (x"4c",x"fb",x"87",x"c2"),
   130 => (x"99",x"c1",x"49",x"73"),
   131 => (x"c3",x"87",x"cd",x"05"),
   132 => (x"c4",x"e0",x"49",x"f4"),
   133 => (x"c2",x"49",x"70",x"87"),
   134 => (x"87",x"c2",x"02",x"99"),
   135 => (x"49",x"73",x"4c",x"fa"),
   136 => (x"ce",x"05",x"99",x"c8"),
   137 => (x"49",x"f5",x"c3",x"87"),
   138 => (x"87",x"ed",x"df",x"ff"),
   139 => (x"99",x"c2",x"49",x"70"),
   140 => (x"c2",x"87",x"d5",x"02"),
   141 => (x"02",x"bf",x"d2",x"ee"),
   142 => (x"c1",x"48",x"87",x"ca"),
   143 => (x"d6",x"ee",x"c2",x"88"),
   144 => (x"87",x"c2",x"c0",x"58"),
   145 => (x"4d",x"c1",x"4c",x"ff"),
   146 => (x"99",x"c4",x"49",x"73"),
   147 => (x"c3",x"87",x"ce",x"05"),
   148 => (x"df",x"ff",x"49",x"f2"),
   149 => (x"49",x"70",x"87",x"c3"),
   150 => (x"dc",x"02",x"99",x"c2"),
   151 => (x"d2",x"ee",x"c2",x"87"),
   152 => (x"c7",x"48",x"7e",x"bf"),
   153 => (x"c0",x"03",x"a8",x"b7"),
   154 => (x"48",x"6e",x"87",x"cb"),
   155 => (x"ee",x"c2",x"80",x"c1"),
   156 => (x"c2",x"c0",x"58",x"d6"),
   157 => (x"c1",x"4c",x"fe",x"87"),
   158 => (x"49",x"fd",x"c3",x"4d"),
   159 => (x"87",x"d9",x"de",x"ff"),
   160 => (x"99",x"c2",x"49",x"70"),
   161 => (x"87",x"d5",x"c0",x"02"),
   162 => (x"bf",x"d2",x"ee",x"c2"),
   163 => (x"87",x"c9",x"c0",x"02"),
   164 => (x"48",x"d2",x"ee",x"c2"),
   165 => (x"c2",x"c0",x"78",x"c0"),
   166 => (x"c1",x"4c",x"fd",x"87"),
   167 => (x"49",x"fa",x"c3",x"4d"),
   168 => (x"87",x"f5",x"dd",x"ff"),
   169 => (x"99",x"c2",x"49",x"70"),
   170 => (x"87",x"d9",x"c0",x"02"),
   171 => (x"bf",x"d2",x"ee",x"c2"),
   172 => (x"a8",x"b7",x"c7",x"48"),
   173 => (x"87",x"c9",x"c0",x"03"),
   174 => (x"48",x"d2",x"ee",x"c2"),
   175 => (x"c2",x"c0",x"78",x"c7"),
   176 => (x"c1",x"4c",x"fc",x"87"),
   177 => (x"ac",x"b7",x"c0",x"4d"),
   178 => (x"87",x"d1",x"c0",x"03"),
   179 => (x"c1",x"4a",x"66",x"c4"),
   180 => (x"02",x"6a",x"82",x"d8"),
   181 => (x"6a",x"87",x"c6",x"c0"),
   182 => (x"73",x"49",x"74",x"4b"),
   183 => (x"c3",x"1e",x"c0",x"0f"),
   184 => (x"da",x"c1",x"1e",x"f0"),
   185 => (x"87",x"e6",x"f6",x"49"),
   186 => (x"98",x"70",x"86",x"c8"),
   187 => (x"87",x"e2",x"c0",x"02"),
   188 => (x"c2",x"48",x"a6",x"c8"),
   189 => (x"78",x"bf",x"d2",x"ee"),
   190 => (x"cb",x"49",x"66",x"c8"),
   191 => (x"48",x"66",x"c4",x"91"),
   192 => (x"7e",x"70",x"80",x"71"),
   193 => (x"c0",x"02",x"bf",x"6e"),
   194 => (x"bf",x"6e",x"87",x"c8"),
   195 => (x"49",x"66",x"c8",x"4b"),
   196 => (x"9d",x"75",x"0f",x"73"),
   197 => (x"87",x"c8",x"c0",x"02"),
   198 => (x"bf",x"d2",x"ee",x"c2"),
   199 => (x"87",x"d4",x"f2",x"49"),
   200 => (x"bf",x"f4",x"ce",x"c2"),
   201 => (x"87",x"dd",x"c0",x"02"),
   202 => (x"87",x"d8",x"c2",x"49"),
   203 => (x"c0",x"02",x"98",x"70"),
   204 => (x"ee",x"c2",x"87",x"d3"),
   205 => (x"f1",x"49",x"bf",x"d2"),
   206 => (x"49",x"c0",x"87",x"fa"),
   207 => (x"c2",x"87",x"da",x"f3"),
   208 => (x"c0",x"48",x"f4",x"ce"),
   209 => (x"f2",x"8e",x"f4",x"78"),
   210 => (x"5e",x"0e",x"87",x"f4"),
   211 => (x"0e",x"5d",x"5c",x"5b"),
   212 => (x"c2",x"4c",x"71",x"1e"),
   213 => (x"49",x"bf",x"ce",x"ee"),
   214 => (x"4d",x"a1",x"cd",x"c1"),
   215 => (x"69",x"81",x"d1",x"c1"),
   216 => (x"02",x"9c",x"74",x"7e"),
   217 => (x"a5",x"c4",x"87",x"cf"),
   218 => (x"c2",x"7b",x"74",x"4b"),
   219 => (x"49",x"bf",x"ce",x"ee"),
   220 => (x"6e",x"87",x"d3",x"f2"),
   221 => (x"05",x"9c",x"74",x"7b"),
   222 => (x"4b",x"c0",x"87",x"c4"),
   223 => (x"4b",x"c1",x"87",x"c2"),
   224 => (x"d4",x"f2",x"49",x"73"),
   225 => (x"02",x"66",x"d4",x"87"),
   226 => (x"c0",x"49",x"87",x"c8"),
   227 => (x"4a",x"70",x"87",x"ea"),
   228 => (x"4a",x"c0",x"87",x"c2"),
   229 => (x"5a",x"f8",x"ce",x"c2"),
   230 => (x"87",x"e2",x"f1",x"26"),
   231 => (x"14",x"11",x"12",x"58"),
   232 => (x"23",x"1c",x"1b",x"1d"),
   233 => (x"94",x"91",x"59",x"5a"),
   234 => (x"f4",x"eb",x"f2",x"f5"),
   235 => (x"00",x"00",x"00",x"00"),
   236 => (x"00",x"00",x"00",x"00"),
   237 => (x"00",x"00",x"00",x"00"),
   238 => (x"ff",x"4a",x"71",x"1e"),
   239 => (x"72",x"49",x"bf",x"c8"),
   240 => (x"4f",x"26",x"48",x"a1"),
   241 => (x"bf",x"c8",x"ff",x"1e"),
   242 => (x"c0",x"c0",x"fe",x"89"),
   243 => (x"a9",x"c0",x"c0",x"c0"),
   244 => (x"c0",x"87",x"c4",x"01"),
   245 => (x"c1",x"87",x"c2",x"4a"),
   246 => (x"26",x"48",x"72",x"4a"),
   247 => (x"5b",x"5e",x"0e",x"4f"),
   248 => (x"71",x"0e",x"5d",x"5c"),
   249 => (x"4c",x"d4",x"ff",x"4b"),
   250 => (x"c0",x"48",x"66",x"d0"),
   251 => (x"ff",x"49",x"d6",x"78"),
   252 => (x"c3",x"87",x"e6",x"da"),
   253 => (x"49",x"6c",x"7c",x"ff"),
   254 => (x"71",x"99",x"ff",x"c3"),
   255 => (x"f0",x"c3",x"49",x"4d"),
   256 => (x"a9",x"e0",x"c1",x"99"),
   257 => (x"c3",x"87",x"cb",x"05"),
   258 => (x"48",x"6c",x"7c",x"ff"),
   259 => (x"66",x"d0",x"98",x"c3"),
   260 => (x"ff",x"c3",x"78",x"08"),
   261 => (x"49",x"4a",x"6c",x"7c"),
   262 => (x"ff",x"c3",x"31",x"c8"),
   263 => (x"71",x"4a",x"6c",x"7c"),
   264 => (x"c8",x"49",x"72",x"b2"),
   265 => (x"7c",x"ff",x"c3",x"31"),
   266 => (x"b2",x"71",x"4a",x"6c"),
   267 => (x"31",x"c8",x"49",x"72"),
   268 => (x"6c",x"7c",x"ff",x"c3"),
   269 => (x"ff",x"b2",x"71",x"4a"),
   270 => (x"e0",x"c0",x"48",x"d0"),
   271 => (x"02",x"9b",x"73",x"78"),
   272 => (x"7b",x"72",x"87",x"c2"),
   273 => (x"4d",x"26",x"48",x"75"),
   274 => (x"4b",x"26",x"4c",x"26"),
   275 => (x"26",x"1e",x"4f",x"26"),
   276 => (x"5b",x"5e",x"0e",x"4f"),
   277 => (x"86",x"f8",x"0e",x"5c"),
   278 => (x"a6",x"c8",x"1e",x"76"),
   279 => (x"87",x"fd",x"fd",x"49"),
   280 => (x"4b",x"70",x"86",x"c4"),
   281 => (x"a8",x"c2",x"48",x"6e"),
   282 => (x"87",x"f0",x"c2",x"03"),
   283 => (x"f0",x"c3",x"4a",x"73"),
   284 => (x"aa",x"d0",x"c1",x"9a"),
   285 => (x"c1",x"87",x"c7",x"02"),
   286 => (x"c2",x"05",x"aa",x"e0"),
   287 => (x"49",x"73",x"87",x"de"),
   288 => (x"c3",x"02",x"99",x"c8"),
   289 => (x"87",x"c6",x"ff",x"87"),
   290 => (x"9c",x"c3",x"4c",x"73"),
   291 => (x"c1",x"05",x"ac",x"c2"),
   292 => (x"66",x"c4",x"87",x"c2"),
   293 => (x"71",x"31",x"c9",x"49"),
   294 => (x"4a",x"66",x"c4",x"1e"),
   295 => (x"ee",x"c2",x"92",x"d4"),
   296 => (x"81",x"72",x"49",x"d6"),
   297 => (x"87",x"c7",x"d4",x"fe"),
   298 => (x"d7",x"ff",x"49",x"d8"),
   299 => (x"c0",x"c8",x"87",x"eb"),
   300 => (x"c6",x"dd",x"c2",x"1e"),
   301 => (x"e2",x"f0",x"fd",x"49"),
   302 => (x"48",x"d0",x"ff",x"87"),
   303 => (x"c2",x"78",x"e0",x"c0"),
   304 => (x"cc",x"1e",x"c6",x"dd"),
   305 => (x"92",x"d4",x"4a",x"66"),
   306 => (x"49",x"d6",x"ee",x"c2"),
   307 => (x"d2",x"fe",x"81",x"72"),
   308 => (x"86",x"cc",x"87",x"da"),
   309 => (x"c1",x"05",x"ac",x"c1"),
   310 => (x"66",x"c4",x"87",x"c2"),
   311 => (x"71",x"31",x"c9",x"49"),
   312 => (x"4a",x"66",x"c4",x"1e"),
   313 => (x"ee",x"c2",x"92",x"d4"),
   314 => (x"81",x"72",x"49",x"d6"),
   315 => (x"87",x"ff",x"d2",x"fe"),
   316 => (x"1e",x"c6",x"dd",x"c2"),
   317 => (x"d4",x"4a",x"66",x"c8"),
   318 => (x"d6",x"ee",x"c2",x"92"),
   319 => (x"fe",x"81",x"72",x"49"),
   320 => (x"d7",x"87",x"e6",x"d0"),
   321 => (x"d0",x"d6",x"ff",x"49"),
   322 => (x"1e",x"c0",x"c8",x"87"),
   323 => (x"49",x"c6",x"dd",x"c2"),
   324 => (x"87",x"f1",x"ee",x"fd"),
   325 => (x"d0",x"ff",x"86",x"cc"),
   326 => (x"78",x"e0",x"c0",x"48"),
   327 => (x"e7",x"fc",x"8e",x"f8"),
   328 => (x"5b",x"5e",x"0e",x"87"),
   329 => (x"1e",x"0e",x"5d",x"5c"),
   330 => (x"d4",x"ff",x"4d",x"71"),
   331 => (x"7e",x"66",x"d4",x"4c"),
   332 => (x"a8",x"b7",x"c3",x"48"),
   333 => (x"c0",x"87",x"c5",x"06"),
   334 => (x"87",x"e2",x"c1",x"48"),
   335 => (x"e0",x"fe",x"49",x"75"),
   336 => (x"1e",x"75",x"87",x"fe"),
   337 => (x"d4",x"4b",x"66",x"c4"),
   338 => (x"d6",x"ee",x"c2",x"93"),
   339 => (x"fe",x"49",x"73",x"83"),
   340 => (x"c8",x"87",x"fa",x"cb"),
   341 => (x"ff",x"4b",x"6b",x"83"),
   342 => (x"e1",x"c8",x"48",x"d0"),
   343 => (x"73",x"7c",x"dd",x"78"),
   344 => (x"99",x"ff",x"c3",x"49"),
   345 => (x"49",x"73",x"7c",x"71"),
   346 => (x"c3",x"29",x"b7",x"c8"),
   347 => (x"7c",x"71",x"99",x"ff"),
   348 => (x"b7",x"d0",x"49",x"73"),
   349 => (x"99",x"ff",x"c3",x"29"),
   350 => (x"49",x"73",x"7c",x"71"),
   351 => (x"71",x"29",x"b7",x"d8"),
   352 => (x"7c",x"7c",x"c0",x"7c"),
   353 => (x"7c",x"7c",x"7c",x"7c"),
   354 => (x"7c",x"7c",x"7c",x"7c"),
   355 => (x"e0",x"c0",x"7c",x"7c"),
   356 => (x"1e",x"66",x"c4",x"78"),
   357 => (x"d4",x"ff",x"49",x"dc"),
   358 => (x"86",x"c8",x"87",x"e4"),
   359 => (x"fa",x"26",x"48",x"73"),
   360 => (x"5e",x"0e",x"87",x"e4"),
   361 => (x"0e",x"5d",x"5c",x"5b"),
   362 => (x"ff",x"7e",x"71",x"1e"),
   363 => (x"1e",x"6e",x"4b",x"d4"),
   364 => (x"49",x"fe",x"ee",x"c2"),
   365 => (x"87",x"d5",x"ca",x"fe"),
   366 => (x"4d",x"70",x"86",x"c4"),
   367 => (x"c3",x"c3",x"02",x"9d"),
   368 => (x"c6",x"ef",x"c2",x"87"),
   369 => (x"49",x"6e",x"4c",x"bf"),
   370 => (x"87",x"f4",x"de",x"fe"),
   371 => (x"c8",x"48",x"d0",x"ff"),
   372 => (x"d6",x"c1",x"78",x"c5"),
   373 => (x"15",x"4a",x"c0",x"7b"),
   374 => (x"c0",x"82",x"c1",x"7b"),
   375 => (x"04",x"aa",x"b7",x"e0"),
   376 => (x"d0",x"ff",x"87",x"f5"),
   377 => (x"c8",x"78",x"c4",x"48"),
   378 => (x"d3",x"c1",x"78",x"c5"),
   379 => (x"c4",x"7b",x"c1",x"7b"),
   380 => (x"02",x"9c",x"74",x"78"),
   381 => (x"c2",x"87",x"fc",x"c1"),
   382 => (x"c8",x"7e",x"c6",x"dd"),
   383 => (x"c0",x"8c",x"4d",x"c0"),
   384 => (x"c6",x"03",x"ac",x"b7"),
   385 => (x"a4",x"c0",x"c8",x"87"),
   386 => (x"c2",x"4c",x"c0",x"4d"),
   387 => (x"bf",x"97",x"f7",x"e9"),
   388 => (x"02",x"99",x"d0",x"49"),
   389 => (x"1e",x"c0",x"87",x"d2"),
   390 => (x"49",x"fe",x"ee",x"c2"),
   391 => (x"87",x"c9",x"cc",x"fe"),
   392 => (x"49",x"70",x"86",x"c4"),
   393 => (x"87",x"ef",x"c0",x"4a"),
   394 => (x"1e",x"c6",x"dd",x"c2"),
   395 => (x"49",x"fe",x"ee",x"c2"),
   396 => (x"87",x"f5",x"cb",x"fe"),
   397 => (x"49",x"70",x"86",x"c4"),
   398 => (x"48",x"d0",x"ff",x"4a"),
   399 => (x"c1",x"78",x"c5",x"c8"),
   400 => (x"97",x"6e",x"7b",x"d4"),
   401 => (x"48",x"6e",x"7b",x"bf"),
   402 => (x"7e",x"70",x"80",x"c1"),
   403 => (x"ff",x"05",x"8d",x"c1"),
   404 => (x"d0",x"ff",x"87",x"f0"),
   405 => (x"72",x"78",x"c4",x"48"),
   406 => (x"87",x"c5",x"05",x"9a"),
   407 => (x"e5",x"c0",x"48",x"c0"),
   408 => (x"c2",x"1e",x"c1",x"87"),
   409 => (x"fe",x"49",x"fe",x"ee"),
   410 => (x"c4",x"87",x"dd",x"c9"),
   411 => (x"05",x"9c",x"74",x"86"),
   412 => (x"ff",x"87",x"c4",x"fe"),
   413 => (x"c5",x"c8",x"48",x"d0"),
   414 => (x"7b",x"d3",x"c1",x"78"),
   415 => (x"78",x"c4",x"7b",x"c0"),
   416 => (x"87",x"c2",x"48",x"c1"),
   417 => (x"26",x"26",x"48",x"c0"),
   418 => (x"26",x"4c",x"26",x"4d"),
   419 => (x"0e",x"4f",x"26",x"4b"),
   420 => (x"0e",x"5c",x"5b",x"5e"),
   421 => (x"66",x"cc",x"4b",x"71"),
   422 => (x"4c",x"87",x"d8",x"02"),
   423 => (x"02",x"8c",x"f0",x"c0"),
   424 => (x"4a",x"74",x"87",x"d8"),
   425 => (x"d1",x"02",x"8a",x"c1"),
   426 => (x"cd",x"02",x"8a",x"87"),
   427 => (x"c9",x"02",x"8a",x"87"),
   428 => (x"73",x"87",x"d7",x"87"),
   429 => (x"87",x"ea",x"fb",x"49"),
   430 => (x"1e",x"74",x"87",x"d0"),
   431 => (x"e0",x"f9",x"49",x"c0"),
   432 => (x"73",x"1e",x"74",x"87"),
   433 => (x"87",x"d9",x"f9",x"49"),
   434 => (x"fc",x"fe",x"86",x"c8"),
   435 => (x"c2",x"1e",x"00",x"87"),
   436 => (x"49",x"bf",x"dc",x"dc"),
   437 => (x"dc",x"c2",x"b9",x"c1"),
   438 => (x"d4",x"ff",x"59",x"e0"),
   439 => (x"78",x"ff",x"c3",x"48"),
   440 => (x"c8",x"48",x"d0",x"ff"),
   441 => (x"d4",x"ff",x"78",x"e1"),
   442 => (x"c4",x"78",x"c1",x"48"),
   443 => (x"ff",x"78",x"71",x"31"),
   444 => (x"e0",x"c0",x"48",x"d0"),
   445 => (x"1e",x"4f",x"26",x"78"),
   446 => (x"1e",x"d0",x"dc",x"c2"),
   447 => (x"49",x"fe",x"ee",x"c2"),
   448 => (x"87",x"c9",x"c5",x"fe"),
   449 => (x"98",x"70",x"86",x"c4"),
   450 => (x"ff",x"87",x"c3",x"02"),
   451 => (x"4f",x"26",x"87",x"c0"),
   452 => (x"48",x"4b",x"35",x"31"),
   453 => (x"20",x"20",x"20",x"5a"),
   454 => (x"00",x"47",x"46",x"43"),
   455 => (x"00",x"00",x"00",x"00"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

