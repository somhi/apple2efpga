/home/jordi/FPGAs/FPGA-Deca/Deca_17/_A_GITHUB/Apple2efpga_dmty_cape/Apple2efpga_dmty_3p_cape/demistify/xilinx/keyboard.vhd